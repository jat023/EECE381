// nios_system.v

// Generated using ACDS version 13.0sp1 232 at 2015.04.08.11:25:48

`timescale 1 ps / 1 ps
module nios_system (
		input  wire        clk_clk,                     //              clk.clk
		input  wire [3:0]  keys_export,                 //             keys.export
		output wire [3:0]  leds_export,                 //             leds.export
		input  wire        reset_reset_n,               //            reset.reset_n
		output wire [11:0] sdram_wire_addr,             //       sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,               //                 .ba
		output wire        sdram_wire_cas_n,            //                 .cas_n
		output wire        sdram_wire_cke,              //                 .cke
		output wire        sdram_wire_cs_n,             //                 .cs_n
		inout  wire [15:0] sdram_wire_dq,               //                 .dq
		output wire [1:0]  sdram_wire_dqm,              //                 .dqm
		output wire        sdram_wire_ras_n,            //                 .ras_n
		output wire        sdram_wire_we_n,             //                 .we_n
		output wire        sdram_clk_clk,               //        sdram_clk.clk
		inout  wire [7:0]  lcd_data_DATA,               //         lcd_data.DATA
		output wire        lcd_data_ON,                 //                 .ON
		output wire        lcd_data_BLON,               //                 .BLON
		output wire        lcd_data_EN,                 //                 .EN
		output wire        lcd_data_RS,                 //                 .RS
		output wire        lcd_data_RW,                 //                 .RW
		inout  wire        sd_card_b_SD_cmd,            //          sd_card.b_SD_cmd
		inout  wire        sd_card_b_SD_dat,            //                 .b_SD_dat
		inout  wire        sd_card_b_SD_dat3,           //                 .b_SD_dat3
		output wire        sd_card_o_SD_clock,          //                 .o_SD_clock
		output wire        audio_clk_clk,               //        audio_clk.clk
		input  wire        clk_27_clk,                  //           clk_27.clk
		inout  wire [15:0] sram_pixel_DQ,               //       sram_pixel.DQ
		output wire [17:0] sram_pixel_ADDR,             //                 .ADDR
		output wire        sram_pixel_LB_N,             //                 .LB_N
		output wire        sram_pixel_UB_N,             //                 .UB_N
		output wire        sram_pixel_CE_N,             //                 .CE_N
		output wire        sram_pixel_OE_N,             //                 .OE_N
		output wire        sram_pixel_WE_N,             //                 .WE_N
		output wire        vga_controller_CLK,          //   vga_controller.CLK
		output wire        vga_controller_HS,           //                 .HS
		output wire        vga_controller_VS,           //                 .VS
		output wire        vga_controller_BLANK,        //                 .BLANK
		output wire        vga_controller_SYNC,         //                 .SYNC
		output wire [9:0]  vga_controller_R,            //                 .R
		output wire [9:0]  vga_controller_G,            //                 .G
		output wire [9:0]  vga_controller_B,            //                 .B
		input  wire [11:0] dual_port_ram_s2_address,    // dual_port_ram_s2.address
		input  wire        dual_port_ram_s2_chipselect, //                 .chipselect
		input  wire        dual_port_ram_s2_clken,      //                 .clken
		input  wire        dual_port_ram_s2_write,      //                 .write
		output wire [7:0]  dual_port_ram_s2_readdata,   //                 .readdata
		input  wire [7:0]  dual_port_ram_s2_writedata,  //                 .writedata
		input  wire        clk_pi_clk,                  //           clk_pi.clk
		output wire        de2_ack_export,              //          de2_ack.export
		input  wire        pi_request_export            //       pi_request.export
	);

	wire          clocks_sys_clk_clk;                                                                                         // clocks:sys_clk -> [LEDs:clk, LEDs_s1_translator:clk, LEDs_s1_translator_avalon_universal_slave_0_agent:clk, LEDs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, addr_router:clk, addr_router_001:clk, addr_router_002:clk, addr_router_003:clk, burst_adapter:clk, burst_adapter_001:clk, burst_adapter_002:clk, burst_adapter_003:clk, character_lcd_0:clk, character_lcd_0_avalon_lcd_slave_translator:clk, character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:clk, character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, cmd_xbar_demux:clk, cmd_xbar_demux_001:clk, cmd_xbar_demux_002:clk, cmd_xbar_demux_003:clk, cmd_xbar_mux:clk, cmd_xbar_mux_001:clk, cmd_xbar_mux_002:clk, cmd_xbar_mux_003:clk, cmd_xbar_mux_004:clk, cmd_xbar_mux_005:clk, cmd_xbar_mux_010:clk, de2_ack:clk, de2_ack_s1_translator:clk, de2_ack_s1_translator_avalon_universal_slave_0_agent:clk, de2_ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, dual_port_ram:clk, dual_port_ram_s1_translator:clk, dual_port_ram_s1_translator_avalon_universal_slave_0_agent:clk, dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, id_router:clk, id_router_001:clk, id_router_002:clk, id_router_003:clk, id_router_004:clk, id_router_005:clk, id_router_006:clk, id_router_007:clk, id_router_008:clk, id_router_009:clk, id_router_010:clk, id_router_011:clk, id_router_012:clk, id_router_013:clk, id_router_014:clk, id_router_015:clk, irq_mapper:clk, jtag_uart_0:clk, jtag_uart_0_avalon_jtag_slave_translator:clk, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:clk, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, keys:clk, keys_s1_translator:clk, keys_s1_translator_avalon_universal_slave_0_agent:clk, keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, line_drawer_0:clk, line_drawer_0_avalon_master_translator:clk, line_drawer_0_avalon_master_translator_avalon_universal_master_0_agent:clk, line_drawer_0_avalon_slave_0_translator:clk, line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:clk, line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, nios2_qsys_0:clk, nios2_qsys_0_data_master_translator:clk, nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:clk, nios2_qsys_0_instruction_master_translator:clk, nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:clk, nios2_qsys_0_jtag_debug_module_translator:clk, nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:clk, nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, onchip_memory2_0:clk, onchip_memory2_0_s1_translator:clk, onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:clk, onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pi_request:clk, pi_request_s1_translator:clk, pi_request_s1_translator_avalon_universal_slave_0_agent:clk, pi_request_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pixel_buffer:clk, pixel_buffer_avalon_sram_slave_translator:clk, pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:clk, pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pixel_buffer_dma:clk, pixel_buffer_dma_avalon_control_slave_translator:clk, pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:clk, pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pixel_buffer_dma_avalon_pixel_dma_master_translator:clk, pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:clk, rgb_sampler:clk, rsp_xbar_demux:clk, rsp_xbar_demux_001:clk, rsp_xbar_demux_002:clk, rsp_xbar_demux_003:clk, rsp_xbar_demux_004:clk, rsp_xbar_demux_005:clk, rsp_xbar_demux_006:clk, rsp_xbar_demux_007:clk, rsp_xbar_demux_008:clk, rsp_xbar_demux_009:clk, rsp_xbar_demux_010:clk, rsp_xbar_demux_011:clk, rsp_xbar_demux_012:clk, rsp_xbar_demux_013:clk, rsp_xbar_demux_014:clk, rsp_xbar_demux_015:clk, rsp_xbar_mux:clk, rsp_xbar_mux_001:clk, rst_controller:clk, scaler:clk, sd_card:i_clock, sd_card_avalon_sdcard_slave_translator:clk, sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:clk, sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, sdram:clk, sdram_s1_translator:clk, sdram_s1_translator_avalon_universal_slave_0_agent:clk, sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, timer_system:clk, timer_system_s1_translator:clk, timer_system_s1_translator_avalon_universal_slave_0_agent:clk, timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, timer_timestamp:clk, timer_timestamp_s1_translator:clk, timer_timestamp_s1_translator_avalon_universal_slave_0_agent:clk, timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, video_fifo:clk_stream_in, width_adapter:clk, width_adapter_001:clk, width_adapter_002:clk, width_adapter_003:clk, width_adapter_004:clk, width_adapter_005:clk, width_adapter_006:clk, width_adapter_007:clk, width_adapter_008:clk, width_adapter_009:clk]
	wire          rgb_sampler_avalon_rgb_source_endofpacket;                                                                  // rgb_sampler:stream_out_endofpacket -> scaler:stream_in_endofpacket
	wire          rgb_sampler_avalon_rgb_source_valid;                                                                        // rgb_sampler:stream_out_valid -> scaler:stream_in_valid
	wire          rgb_sampler_avalon_rgb_source_startofpacket;                                                                // rgb_sampler:stream_out_startofpacket -> scaler:stream_in_startofpacket
	wire   [29:0] rgb_sampler_avalon_rgb_source_data;                                                                         // rgb_sampler:stream_out_data -> scaler:stream_in_data
	wire          rgb_sampler_avalon_rgb_source_ready;                                                                        // scaler:stream_in_ready -> rgb_sampler:stream_out_ready
	wire          clocks_vga_clk_clk;                                                                                         // clocks:VGA_CLK -> [rst_controller_002:clk, vga_controller:clk, video_fifo:clk_stream_out]
	wire          video_fifo_avalon_dc_buffer_source_endofpacket;                                                             // video_fifo:stream_out_endofpacket -> vga_controller:endofpacket
	wire          video_fifo_avalon_dc_buffer_source_valid;                                                                   // video_fifo:stream_out_valid -> vga_controller:valid
	wire          video_fifo_avalon_dc_buffer_source_startofpacket;                                                           // video_fifo:stream_out_startofpacket -> vga_controller:startofpacket
	wire   [29:0] video_fifo_avalon_dc_buffer_source_data;                                                                    // video_fifo:stream_out_data -> vga_controller:data
	wire          video_fifo_avalon_dc_buffer_source_ready;                                                                   // vga_controller:ready -> video_fifo:stream_out_ready
	wire          scaler_avalon_scaler_source_endofpacket;                                                                    // scaler:stream_out_endofpacket -> video_fifo:stream_in_endofpacket
	wire          scaler_avalon_scaler_source_valid;                                                                          // scaler:stream_out_valid -> video_fifo:stream_in_valid
	wire          scaler_avalon_scaler_source_startofpacket;                                                                  // scaler:stream_out_startofpacket -> video_fifo:stream_in_startofpacket
	wire   [29:0] scaler_avalon_scaler_source_data;                                                                           // scaler:stream_out_data -> video_fifo:stream_in_data
	wire          scaler_avalon_scaler_source_ready;                                                                          // video_fifo:stream_in_ready -> scaler:stream_out_ready
	wire          pixel_buffer_dma_avalon_pixel_source_endofpacket;                                                           // pixel_buffer_dma:stream_endofpacket -> rgb_sampler:stream_in_endofpacket
	wire          pixel_buffer_dma_avalon_pixel_source_valid;                                                                 // pixel_buffer_dma:stream_valid -> rgb_sampler:stream_in_valid
	wire          pixel_buffer_dma_avalon_pixel_source_startofpacket;                                                         // pixel_buffer_dma:stream_startofpacket -> rgb_sampler:stream_in_startofpacket
	wire   [15:0] pixel_buffer_dma_avalon_pixel_source_data;                                                                  // pixel_buffer_dma:stream_data -> rgb_sampler:stream_in_data
	wire          pixel_buffer_dma_avalon_pixel_source_ready;                                                                 // rgb_sampler:stream_in_ready -> pixel_buffer_dma:stream_ready
	wire          nios2_qsys_0_instruction_master_waitrequest;                                                                // nios2_qsys_0_instruction_master_translator:av_waitrequest -> nios2_qsys_0:i_waitrequest
	wire   [24:0] nios2_qsys_0_instruction_master_address;                                                                    // nios2_qsys_0:i_address -> nios2_qsys_0_instruction_master_translator:av_address
	wire          nios2_qsys_0_instruction_master_read;                                                                       // nios2_qsys_0:i_read -> nios2_qsys_0_instruction_master_translator:av_read
	wire   [31:0] nios2_qsys_0_instruction_master_readdata;                                                                   // nios2_qsys_0_instruction_master_translator:av_readdata -> nios2_qsys_0:i_readdata
	wire          nios2_qsys_0_data_master_waitrequest;                                                                       // nios2_qsys_0_data_master_translator:av_waitrequest -> nios2_qsys_0:d_waitrequest
	wire   [31:0] nios2_qsys_0_data_master_writedata;                                                                         // nios2_qsys_0:d_writedata -> nios2_qsys_0_data_master_translator:av_writedata
	wire   [24:0] nios2_qsys_0_data_master_address;                                                                           // nios2_qsys_0:d_address -> nios2_qsys_0_data_master_translator:av_address
	wire          nios2_qsys_0_data_master_write;                                                                             // nios2_qsys_0:d_write -> nios2_qsys_0_data_master_translator:av_write
	wire          nios2_qsys_0_data_master_read;                                                                              // nios2_qsys_0:d_read -> nios2_qsys_0_data_master_translator:av_read
	wire   [31:0] nios2_qsys_0_data_master_readdata;                                                                          // nios2_qsys_0_data_master_translator:av_readdata -> nios2_qsys_0:d_readdata
	wire          nios2_qsys_0_data_master_debugaccess;                                                                       // nios2_qsys_0:jtag_debug_module_debugaccess_to_roms -> nios2_qsys_0_data_master_translator:av_debugaccess
	wire    [3:0] nios2_qsys_0_data_master_byteenable;                                                                        // nios2_qsys_0:d_byteenable -> nios2_qsys_0_data_master_translator:av_byteenable
	wire          pixel_buffer_dma_avalon_pixel_dma_master_waitrequest;                                                       // pixel_buffer_dma_avalon_pixel_dma_master_translator:av_waitrequest -> pixel_buffer_dma:master_waitrequest
	wire   [31:0] pixel_buffer_dma_avalon_pixel_dma_master_address;                                                           // pixel_buffer_dma:master_address -> pixel_buffer_dma_avalon_pixel_dma_master_translator:av_address
	wire          pixel_buffer_dma_avalon_pixel_dma_master_lock;                                                              // pixel_buffer_dma:master_arbiterlock -> pixel_buffer_dma_avalon_pixel_dma_master_translator:av_lock
	wire          pixel_buffer_dma_avalon_pixel_dma_master_read;                                                              // pixel_buffer_dma:master_read -> pixel_buffer_dma_avalon_pixel_dma_master_translator:av_read
	wire   [15:0] pixel_buffer_dma_avalon_pixel_dma_master_readdata;                                                          // pixel_buffer_dma_avalon_pixel_dma_master_translator:av_readdata -> pixel_buffer_dma:master_readdata
	wire          pixel_buffer_dma_avalon_pixel_dma_master_readdatavalid;                                                     // pixel_buffer_dma_avalon_pixel_dma_master_translator:av_readdatavalid -> pixel_buffer_dma:master_readdatavalid
	wire          line_drawer_0_avalon_master_waitrequest;                                                                    // line_drawer_0_avalon_master_translator:av_waitrequest -> line_drawer_0:master_waitrequest
	wire   [31:0] line_drawer_0_avalon_master_address;                                                                        // line_drawer_0:master_addr -> line_drawer_0_avalon_master_translator:av_address
	wire   [15:0] line_drawer_0_avalon_master_writedata;                                                                      // line_drawer_0:master_writedata -> line_drawer_0_avalon_master_translator:av_writedata
	wire          line_drawer_0_avalon_master_write;                                                                          // line_drawer_0:master_wr_en -> line_drawer_0_avalon_master_translator:av_write
	wire          line_drawer_0_avalon_master_read;                                                                           // line_drawer_0:master_rd_en -> line_drawer_0_avalon_master_translator:av_read
	wire   [15:0] line_drawer_0_avalon_master_readdata;                                                                       // line_drawer_0_avalon_master_translator:av_readdata -> line_drawer_0:master_readdata
	wire    [1:0] line_drawer_0_avalon_master_byteenable;                                                                     // line_drawer_0:master_be -> line_drawer_0_avalon_master_translator:av_byteenable
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest;                                  // nios2_qsys_0:jtag_debug_module_waitrequest -> nios2_qsys_0_jtag_debug_module_translator:av_waitrequest
	wire   [31:0] nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                    // nios2_qsys_0_jtag_debug_module_translator:av_writedata -> nios2_qsys_0:jtag_debug_module_writedata
	wire    [8:0] nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_address;                                      // nios2_qsys_0_jtag_debug_module_translator:av_address -> nios2_qsys_0:jtag_debug_module_address
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_write;                                        // nios2_qsys_0_jtag_debug_module_translator:av_write -> nios2_qsys_0:jtag_debug_module_write
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_read;                                         // nios2_qsys_0_jtag_debug_module_translator:av_read -> nios2_qsys_0:jtag_debug_module_read
	wire   [31:0] nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                     // nios2_qsys_0:jtag_debug_module_readdata -> nios2_qsys_0_jtag_debug_module_translator:av_readdata
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                  // nios2_qsys_0_jtag_debug_module_translator:av_debugaccess -> nios2_qsys_0:jtag_debug_module_debugaccess
	wire    [3:0] nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                   // nios2_qsys_0_jtag_debug_module_translator:av_byteenable -> nios2_qsys_0:jtag_debug_module_byteenable
	wire   [31:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_writedata;                                               // onchip_memory2_0_s1_translator:av_writedata -> onchip_memory2_0:writedata
	wire    [9:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_address;                                                 // onchip_memory2_0_s1_translator:av_address -> onchip_memory2_0:address
	wire          onchip_memory2_0_s1_translator_avalon_anti_slave_0_chipselect;                                              // onchip_memory2_0_s1_translator:av_chipselect -> onchip_memory2_0:chipselect
	wire          onchip_memory2_0_s1_translator_avalon_anti_slave_0_clken;                                                   // onchip_memory2_0_s1_translator:av_clken -> onchip_memory2_0:clken
	wire          onchip_memory2_0_s1_translator_avalon_anti_slave_0_write;                                                   // onchip_memory2_0_s1_translator:av_write -> onchip_memory2_0:write
	wire   [31:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_readdata;                                                // onchip_memory2_0:readdata -> onchip_memory2_0_s1_translator:av_readdata
	wire    [3:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_byteenable;                                              // onchip_memory2_0_s1_translator:av_byteenable -> onchip_memory2_0:byteenable
	wire          sdram_s1_translator_avalon_anti_slave_0_waitrequest;                                                        // sdram:za_waitrequest -> sdram_s1_translator:av_waitrequest
	wire   [15:0] sdram_s1_translator_avalon_anti_slave_0_writedata;                                                          // sdram_s1_translator:av_writedata -> sdram:az_data
	wire   [21:0] sdram_s1_translator_avalon_anti_slave_0_address;                                                            // sdram_s1_translator:av_address -> sdram:az_addr
	wire          sdram_s1_translator_avalon_anti_slave_0_chipselect;                                                         // sdram_s1_translator:av_chipselect -> sdram:az_cs
	wire          sdram_s1_translator_avalon_anti_slave_0_write;                                                              // sdram_s1_translator:av_write -> sdram:az_wr_n
	wire          sdram_s1_translator_avalon_anti_slave_0_read;                                                               // sdram_s1_translator:av_read -> sdram:az_rd_n
	wire   [15:0] sdram_s1_translator_avalon_anti_slave_0_readdata;                                                           // sdram:za_data -> sdram_s1_translator:av_readdata
	wire          sdram_s1_translator_avalon_anti_slave_0_readdatavalid;                                                      // sdram:za_valid -> sdram_s1_translator:av_readdatavalid
	wire    [1:0] sdram_s1_translator_avalon_anti_slave_0_byteenable;                                                         // sdram_s1_translator:av_byteenable -> sdram:az_be_n
	wire   [15:0] timer_system_s1_translator_avalon_anti_slave_0_writedata;                                                   // timer_system_s1_translator:av_writedata -> timer_system:writedata
	wire    [2:0] timer_system_s1_translator_avalon_anti_slave_0_address;                                                     // timer_system_s1_translator:av_address -> timer_system:address
	wire          timer_system_s1_translator_avalon_anti_slave_0_chipselect;                                                  // timer_system_s1_translator:av_chipselect -> timer_system:chipselect
	wire          timer_system_s1_translator_avalon_anti_slave_0_write;                                                       // timer_system_s1_translator:av_write -> timer_system:write_n
	wire   [15:0] timer_system_s1_translator_avalon_anti_slave_0_readdata;                                                    // timer_system:readdata -> timer_system_s1_translator:av_readdata
	wire   [15:0] timer_timestamp_s1_translator_avalon_anti_slave_0_writedata;                                                // timer_timestamp_s1_translator:av_writedata -> timer_timestamp:writedata
	wire    [2:0] timer_timestamp_s1_translator_avalon_anti_slave_0_address;                                                  // timer_timestamp_s1_translator:av_address -> timer_timestamp:address
	wire          timer_timestamp_s1_translator_avalon_anti_slave_0_chipselect;                                               // timer_timestamp_s1_translator:av_chipselect -> timer_timestamp:chipselect
	wire          timer_timestamp_s1_translator_avalon_anti_slave_0_write;                                                    // timer_timestamp_s1_translator:av_write -> timer_timestamp:write_n
	wire   [15:0] timer_timestamp_s1_translator_avalon_anti_slave_0_readdata;                                                 // timer_timestamp:readdata -> timer_timestamp_s1_translator:av_readdata
	wire          sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_waitrequest;                                     // sd_card:o_avalon_waitrequest -> sd_card_avalon_sdcard_slave_translator:av_waitrequest
	wire   [31:0] sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_writedata;                                       // sd_card_avalon_sdcard_slave_translator:av_writedata -> sd_card:i_avalon_writedata
	wire    [7:0] sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_address;                                         // sd_card_avalon_sdcard_slave_translator:av_address -> sd_card:i_avalon_address
	wire          sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_chipselect;                                      // sd_card_avalon_sdcard_slave_translator:av_chipselect -> sd_card:i_avalon_chip_select
	wire          sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_write;                                           // sd_card_avalon_sdcard_slave_translator:av_write -> sd_card:i_avalon_write
	wire          sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_read;                                            // sd_card_avalon_sdcard_slave_translator:av_read -> sd_card:i_avalon_read
	wire   [31:0] sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_readdata;                                        // sd_card:o_avalon_readdata -> sd_card_avalon_sdcard_slave_translator:av_readdata
	wire    [3:0] sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_byteenable;                                      // sd_card_avalon_sdcard_slave_translator:av_byteenable -> sd_card:i_avalon_byteenable
	wire    [1:0] keys_s1_translator_avalon_anti_slave_0_address;                                                             // keys_s1_translator:av_address -> keys:address
	wire   [31:0] keys_s1_translator_avalon_anti_slave_0_readdata;                                                            // keys:readdata -> keys_s1_translator:av_readdata
	wire   [31:0] leds_s1_translator_avalon_anti_slave_0_writedata;                                                           // LEDs_s1_translator:av_writedata -> LEDs:writedata
	wire    [1:0] leds_s1_translator_avalon_anti_slave_0_address;                                                             // LEDs_s1_translator:av_address -> LEDs:address
	wire          leds_s1_translator_avalon_anti_slave_0_chipselect;                                                          // LEDs_s1_translator:av_chipselect -> LEDs:chipselect
	wire          leds_s1_translator_avalon_anti_slave_0_write;                                                               // LEDs_s1_translator:av_write -> LEDs:write_n
	wire   [31:0] leds_s1_translator_avalon_anti_slave_0_readdata;                                                            // LEDs:readdata -> LEDs_s1_translator:av_readdata
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                                   // jtag_uart_0:av_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator:av_waitrequest
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                                     // jtag_uart_0_avalon_jtag_slave_translator:av_writedata -> jtag_uart_0:av_writedata
	wire    [0:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                                       // jtag_uart_0_avalon_jtag_slave_translator:av_address -> jtag_uart_0:av_address
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                                    // jtag_uart_0_avalon_jtag_slave_translator:av_chipselect -> jtag_uart_0:av_chipselect
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                         // jtag_uart_0_avalon_jtag_slave_translator:av_write -> jtag_uart_0:av_write_n
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                          // jtag_uart_0_avalon_jtag_slave_translator:av_read -> jtag_uart_0:av_read_n
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                                      // jtag_uart_0:av_readdata -> jtag_uart_0_avalon_jtag_slave_translator:av_readdata
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_waitrequest;                                // character_lcd_0:waitrequest -> character_lcd_0_avalon_lcd_slave_translator:av_waitrequest
	wire    [7:0] character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_writedata;                                  // character_lcd_0_avalon_lcd_slave_translator:av_writedata -> character_lcd_0:writedata
	wire    [0:0] character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_address;                                    // character_lcd_0_avalon_lcd_slave_translator:av_address -> character_lcd_0:address
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_chipselect;                                 // character_lcd_0_avalon_lcd_slave_translator:av_chipselect -> character_lcd_0:chipselect
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_write;                                      // character_lcd_0_avalon_lcd_slave_translator:av_write -> character_lcd_0:write
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_read;                                       // character_lcd_0_avalon_lcd_slave_translator:av_read -> character_lcd_0:read
	wire    [7:0] character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_readdata;                                   // character_lcd_0:readdata -> character_lcd_0_avalon_lcd_slave_translator:av_readdata
	wire   [15:0] pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_writedata;                                    // pixel_buffer_avalon_sram_slave_translator:av_writedata -> pixel_buffer:writedata
	wire   [17:0] pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_address;                                      // pixel_buffer_avalon_sram_slave_translator:av_address -> pixel_buffer:address
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_write;                                        // pixel_buffer_avalon_sram_slave_translator:av_write -> pixel_buffer:write
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_read;                                         // pixel_buffer_avalon_sram_slave_translator:av_read -> pixel_buffer:read
	wire   [15:0] pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_readdata;                                     // pixel_buffer:readdata -> pixel_buffer_avalon_sram_slave_translator:av_readdata
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid;                                // pixel_buffer:readdatavalid -> pixel_buffer_avalon_sram_slave_translator:av_readdatavalid
	wire    [1:0] pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable;                                   // pixel_buffer_avalon_sram_slave_translator:av_byteenable -> pixel_buffer:byteenable
	wire   [31:0] pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_writedata;                             // pixel_buffer_dma_avalon_control_slave_translator:av_writedata -> pixel_buffer_dma:slave_writedata
	wire    [1:0] pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_address;                               // pixel_buffer_dma_avalon_control_slave_translator:av_address -> pixel_buffer_dma:slave_address
	wire          pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_write;                                 // pixel_buffer_dma_avalon_control_slave_translator:av_write -> pixel_buffer_dma:slave_write
	wire          pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_read;                                  // pixel_buffer_dma_avalon_control_slave_translator:av_read -> pixel_buffer_dma:slave_read
	wire   [31:0] pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_readdata;                              // pixel_buffer_dma:slave_readdata -> pixel_buffer_dma_avalon_control_slave_translator:av_readdata
	wire    [3:0] pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_byteenable;                            // pixel_buffer_dma_avalon_control_slave_translator:av_byteenable -> pixel_buffer_dma:slave_byteenable
	wire   [31:0] line_drawer_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata;                                      // line_drawer_0_avalon_slave_0_translator:av_writedata -> line_drawer_0:slave_writedata
	wire    [2:0] line_drawer_0_avalon_slave_0_translator_avalon_anti_slave_0_address;                                        // line_drawer_0_avalon_slave_0_translator:av_address -> line_drawer_0:slave_addr
	wire          line_drawer_0_avalon_slave_0_translator_avalon_anti_slave_0_write;                                          // line_drawer_0_avalon_slave_0_translator:av_write -> line_drawer_0:slave_wr_en
	wire          line_drawer_0_avalon_slave_0_translator_avalon_anti_slave_0_read;                                           // line_drawer_0_avalon_slave_0_translator:av_read -> line_drawer_0:slave_rd_en
	wire   [31:0] line_drawer_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata;                                       // line_drawer_0:slave_readdata -> line_drawer_0_avalon_slave_0_translator:av_readdata
	wire    [7:0] dual_port_ram_s1_translator_avalon_anti_slave_0_writedata;                                                  // dual_port_ram_s1_translator:av_writedata -> dual_port_ram:writedata
	wire   [11:0] dual_port_ram_s1_translator_avalon_anti_slave_0_address;                                                    // dual_port_ram_s1_translator:av_address -> dual_port_ram:address
	wire          dual_port_ram_s1_translator_avalon_anti_slave_0_chipselect;                                                 // dual_port_ram_s1_translator:av_chipselect -> dual_port_ram:chipselect
	wire          dual_port_ram_s1_translator_avalon_anti_slave_0_clken;                                                      // dual_port_ram_s1_translator:av_clken -> dual_port_ram:clken
	wire          dual_port_ram_s1_translator_avalon_anti_slave_0_write;                                                      // dual_port_ram_s1_translator:av_write -> dual_port_ram:write
	wire    [7:0] dual_port_ram_s1_translator_avalon_anti_slave_0_readdata;                                                   // dual_port_ram:readdata -> dual_port_ram_s1_translator:av_readdata
	wire    [1:0] pi_request_s1_translator_avalon_anti_slave_0_address;                                                       // pi_request_s1_translator:av_address -> pi_request:address
	wire   [31:0] pi_request_s1_translator_avalon_anti_slave_0_readdata;                                                      // pi_request:readdata -> pi_request_s1_translator:av_readdata
	wire   [31:0] de2_ack_s1_translator_avalon_anti_slave_0_writedata;                                                        // de2_ack_s1_translator:av_writedata -> de2_ack:writedata
	wire    [1:0] de2_ack_s1_translator_avalon_anti_slave_0_address;                                                          // de2_ack_s1_translator:av_address -> de2_ack:address
	wire          de2_ack_s1_translator_avalon_anti_slave_0_chipselect;                                                       // de2_ack_s1_translator:av_chipselect -> de2_ack:chipselect
	wire          de2_ack_s1_translator_avalon_anti_slave_0_write;                                                            // de2_ack_s1_translator:av_write -> de2_ack:write_n
	wire   [31:0] de2_ack_s1_translator_avalon_anti_slave_0_readdata;                                                         // de2_ack:readdata -> de2_ack_s1_translator:av_readdata
	wire          nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_waitrequest;                           // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_qsys_0_instruction_master_translator:uav_waitrequest
	wire    [2:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_burstcount;                            // nios2_qsys_0_instruction_master_translator:uav_burstcount -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_writedata;                             // nios2_qsys_0_instruction_master_translator:uav_writedata -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_address;                               // nios2_qsys_0_instruction_master_translator:uav_address -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire          nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_lock;                                  // nios2_qsys_0_instruction_master_translator:uav_lock -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire          nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_write;                                 // nios2_qsys_0_instruction_master_translator:uav_write -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire          nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_read;                                  // nios2_qsys_0_instruction_master_translator:uav_read -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdata;                              // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_qsys_0_instruction_master_translator:uav_readdata
	wire          nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_debugaccess;                           // nios2_qsys_0_instruction_master_translator:uav_debugaccess -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_byteenable;                            // nios2_qsys_0_instruction_master_translator:uav_byteenable -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdatavalid;                         // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_qsys_0_instruction_master_translator:uav_readdatavalid
	wire          nios2_qsys_0_data_master_translator_avalon_universal_master_0_waitrequest;                                  // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_qsys_0_data_master_translator:uav_waitrequest
	wire    [2:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_burstcount;                                   // nios2_qsys_0_data_master_translator:uav_burstcount -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_writedata;                                    // nios2_qsys_0_data_master_translator:uav_writedata -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_address;                                      // nios2_qsys_0_data_master_translator:uav_address -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_address
	wire          nios2_qsys_0_data_master_translator_avalon_universal_master_0_lock;                                         // nios2_qsys_0_data_master_translator:uav_lock -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire          nios2_qsys_0_data_master_translator_avalon_universal_master_0_write;                                        // nios2_qsys_0_data_master_translator:uav_write -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_write
	wire          nios2_qsys_0_data_master_translator_avalon_universal_master_0_read;                                         // nios2_qsys_0_data_master_translator:uav_read -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdata;                                     // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_qsys_0_data_master_translator:uav_readdata
	wire          nios2_qsys_0_data_master_translator_avalon_universal_master_0_debugaccess;                                  // nios2_qsys_0_data_master_translator:uav_debugaccess -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_byteenable;                                   // nios2_qsys_0_data_master_translator:uav_byteenable -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdatavalid;                                // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_qsys_0_data_master_translator:uav_readdatavalid
	wire          pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_waitrequest;                  // pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_waitrequest -> pixel_buffer_dma_avalon_pixel_dma_master_translator:uav_waitrequest
	wire    [1:0] pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_burstcount;                   // pixel_buffer_dma_avalon_pixel_dma_master_translator:uav_burstcount -> pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [15:0] pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_writedata;                    // pixel_buffer_dma_avalon_pixel_dma_master_translator:uav_writedata -> pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_address;                      // pixel_buffer_dma_avalon_pixel_dma_master_translator:uav_address -> pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_address
	wire          pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_lock;                         // pixel_buffer_dma_avalon_pixel_dma_master_translator:uav_lock -> pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_lock
	wire          pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_write;                        // pixel_buffer_dma_avalon_pixel_dma_master_translator:uav_write -> pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_write
	wire          pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_read;                         // pixel_buffer_dma_avalon_pixel_dma_master_translator:uav_read -> pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_read
	wire   [15:0] pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdata;                     // pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_readdata -> pixel_buffer_dma_avalon_pixel_dma_master_translator:uav_readdata
	wire          pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_debugaccess;                  // pixel_buffer_dma_avalon_pixel_dma_master_translator:uav_debugaccess -> pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [1:0] pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_byteenable;                   // pixel_buffer_dma_avalon_pixel_dma_master_translator:uav_byteenable -> pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdatavalid;                // pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> pixel_buffer_dma_avalon_pixel_dma_master_translator:uav_readdatavalid
	wire          line_drawer_0_avalon_master_translator_avalon_universal_master_0_waitrequest;                               // line_drawer_0_avalon_master_translator_avalon_universal_master_0_agent:av_waitrequest -> line_drawer_0_avalon_master_translator:uav_waitrequest
	wire    [1:0] line_drawer_0_avalon_master_translator_avalon_universal_master_0_burstcount;                                // line_drawer_0_avalon_master_translator:uav_burstcount -> line_drawer_0_avalon_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [15:0] line_drawer_0_avalon_master_translator_avalon_universal_master_0_writedata;                                 // line_drawer_0_avalon_master_translator:uav_writedata -> line_drawer_0_avalon_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] line_drawer_0_avalon_master_translator_avalon_universal_master_0_address;                                   // line_drawer_0_avalon_master_translator:uav_address -> line_drawer_0_avalon_master_translator_avalon_universal_master_0_agent:av_address
	wire          line_drawer_0_avalon_master_translator_avalon_universal_master_0_lock;                                      // line_drawer_0_avalon_master_translator:uav_lock -> line_drawer_0_avalon_master_translator_avalon_universal_master_0_agent:av_lock
	wire          line_drawer_0_avalon_master_translator_avalon_universal_master_0_write;                                     // line_drawer_0_avalon_master_translator:uav_write -> line_drawer_0_avalon_master_translator_avalon_universal_master_0_agent:av_write
	wire          line_drawer_0_avalon_master_translator_avalon_universal_master_0_read;                                      // line_drawer_0_avalon_master_translator:uav_read -> line_drawer_0_avalon_master_translator_avalon_universal_master_0_agent:av_read
	wire   [15:0] line_drawer_0_avalon_master_translator_avalon_universal_master_0_readdata;                                  // line_drawer_0_avalon_master_translator_avalon_universal_master_0_agent:av_readdata -> line_drawer_0_avalon_master_translator:uav_readdata
	wire          line_drawer_0_avalon_master_translator_avalon_universal_master_0_debugaccess;                               // line_drawer_0_avalon_master_translator:uav_debugaccess -> line_drawer_0_avalon_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [1:0] line_drawer_0_avalon_master_translator_avalon_universal_master_0_byteenable;                                // line_drawer_0_avalon_master_translator:uav_byteenable -> line_drawer_0_avalon_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          line_drawer_0_avalon_master_translator_avalon_universal_master_0_readdatavalid;                             // line_drawer_0_avalon_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> line_drawer_0_avalon_master_translator:uav_readdatavalid
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                    // nios2_qsys_0_jtag_debug_module_translator:uav_waitrequest -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                     // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> nios2_qsys_0_jtag_debug_module_translator:uav_burstcount
	wire   [31:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                      // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> nios2_qsys_0_jtag_debug_module_translator:uav_writedata
	wire   [31:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                        // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> nios2_qsys_0_jtag_debug_module_translator:uav_address
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                          // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> nios2_qsys_0_jtag_debug_module_translator:uav_write
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                           // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> nios2_qsys_0_jtag_debug_module_translator:uav_lock
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                           // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> nios2_qsys_0_jtag_debug_module_translator:uav_read
	wire   [31:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                       // nios2_qsys_0_jtag_debug_module_translator:uav_readdata -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                  // nios2_qsys_0_jtag_debug_module_translator:uav_readdatavalid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                    // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> nios2_qsys_0_jtag_debug_module_translator:uav_debugaccess
	wire    [3:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                     // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> nios2_qsys_0_jtag_debug_module_translator:uav_byteenable
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;             // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                   // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;           // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                    // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                   // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;          // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;        // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                 // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;              // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;               // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;              // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // onchip_memory2_0_s1_translator:uav_waitrequest -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> onchip_memory2_0_s1_translator:uav_burstcount
	wire   [31:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> onchip_memory2_0_s1_translator:uav_writedata
	wire   [31:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                   // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> onchip_memory2_0_s1_translator:uav_address
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                     // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> onchip_memory2_0_s1_translator:uav_write
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                      // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> onchip_memory2_0_s1_translator:uav_lock
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                      // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> onchip_memory2_0_s1_translator:uav_read
	wire   [31:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // onchip_memory2_0_s1_translator:uav_readdata -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // onchip_memory2_0_s1_translator:uav_readdatavalid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> onchip_memory2_0_s1_translator:uav_debugaccess
	wire    [3:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> onchip_memory2_0_s1_translator:uav_byteenable
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                               // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                          // sdram_s1_translator:uav_waitrequest -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [1:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                           // sdram_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sdram_s1_translator:uav_burstcount
	wire   [15:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                            // sdram_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sdram_s1_translator:uav_writedata
	wire   [31:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_address;                                              // sdram_s1_translator_avalon_universal_slave_0_agent:m0_address -> sdram_s1_translator:uav_address
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                // sdram_s1_translator_avalon_universal_slave_0_agent:m0_write -> sdram_s1_translator:uav_write
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                 // sdram_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sdram_s1_translator:uav_lock
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                 // sdram_s1_translator_avalon_universal_slave_0_agent:m0_read -> sdram_s1_translator:uav_read
	wire   [15:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                             // sdram_s1_translator:uav_readdata -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                        // sdram_s1_translator:uav_readdatavalid -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                          // sdram_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sdram_s1_translator:uav_debugaccess
	wire    [1:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                           // sdram_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sdram_s1_translator:uav_byteenable
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                   // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                         // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                 // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [89:0] sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                          // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                         // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                      // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                              // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [89:0] sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                       // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                      // sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                    // sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [17:0] sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                     // sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                    // sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                                    // sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [17:0] sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                                     // sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                                    // sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          timer_system_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                   // timer_system_s1_translator:uav_waitrequest -> timer_system_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] timer_system_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                    // timer_system_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_system_s1_translator:uav_burstcount
	wire   [31:0] timer_system_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                     // timer_system_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_system_s1_translator:uav_writedata
	wire   [31:0] timer_system_s1_translator_avalon_universal_slave_0_agent_m0_address;                                       // timer_system_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_system_s1_translator:uav_address
	wire          timer_system_s1_translator_avalon_universal_slave_0_agent_m0_write;                                         // timer_system_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_system_s1_translator:uav_write
	wire          timer_system_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                          // timer_system_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_system_s1_translator:uav_lock
	wire          timer_system_s1_translator_avalon_universal_slave_0_agent_m0_read;                                          // timer_system_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_system_s1_translator:uav_read
	wire   [31:0] timer_system_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                      // timer_system_s1_translator:uav_readdata -> timer_system_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          timer_system_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                 // timer_system_s1_translator:uav_readdatavalid -> timer_system_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          timer_system_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                   // timer_system_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_system_s1_translator:uav_debugaccess
	wire    [3:0] timer_system_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                    // timer_system_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_system_s1_translator:uav_byteenable
	wire          timer_system_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                            // timer_system_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          timer_system_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                  // timer_system_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          timer_system_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                          // timer_system_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] timer_system_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                   // timer_system_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          timer_system_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                  // timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_system_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                         // timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_system_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                               // timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_system_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                       // timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_system_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                // timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_system_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                               // timer_system_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          timer_system_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                             // timer_system_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_system_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] timer_system_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                              // timer_system_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_system_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          timer_system_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                             // timer_system_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_system_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // timer_timestamp_s1_translator:uav_waitrequest -> timer_timestamp_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // timer_timestamp_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_timestamp_s1_translator:uav_burstcount
	wire   [31:0] timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // timer_timestamp_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_timestamp_s1_translator:uav_writedata
	wire   [31:0] timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_address;                                    // timer_timestamp_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_timestamp_s1_translator:uav_address
	wire          timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_write;                                      // timer_timestamp_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_timestamp_s1_translator:uav_write
	wire          timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                       // timer_timestamp_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_timestamp_s1_translator:uav_lock
	wire          timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_read;                                       // timer_timestamp_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_timestamp_s1_translator:uav_read
	wire   [31:0] timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // timer_timestamp_s1_translator:uav_readdata -> timer_timestamp_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // timer_timestamp_s1_translator:uav_readdatavalid -> timer_timestamp_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // timer_timestamp_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_timestamp_s1_translator:uav_debugaccess
	wire    [3:0] timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // timer_timestamp_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_timestamp_s1_translator:uav_byteenable
	wire          timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // timer_timestamp_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // timer_timestamp_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // timer_timestamp_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                // timer_timestamp_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_timestamp_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_timestamp_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_timestamp_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_timestamp_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_timestamp_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // timer_timestamp_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // timer_timestamp_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_timestamp_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // timer_timestamp_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_timestamp_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // timer_timestamp_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_timestamp_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                       // sd_card_avalon_sdcard_slave_translator:uav_waitrequest -> sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                        // sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sd_card_avalon_sdcard_slave_translator:uav_burstcount
	wire   [31:0] sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                         // sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sd_card_avalon_sdcard_slave_translator:uav_writedata
	wire   [31:0] sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_address;                           // sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_address -> sd_card_avalon_sdcard_slave_translator:uav_address
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_write;                             // sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_write -> sd_card_avalon_sdcard_slave_translator:uav_write
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_lock;                              // sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sd_card_avalon_sdcard_slave_translator:uav_lock
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_read;                              // sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_read -> sd_card_avalon_sdcard_slave_translator:uav_read
	wire   [31:0] sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                          // sd_card_avalon_sdcard_slave_translator:uav_readdata -> sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                     // sd_card_avalon_sdcard_slave_translator:uav_readdatavalid -> sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                       // sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sd_card_avalon_sdcard_slave_translator:uav_debugaccess
	wire    [3:0] sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                        // sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sd_card_avalon_sdcard_slave_translator:uav_byteenable
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                // sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                      // sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;              // sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                       // sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                      // sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;             // sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                   // sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;           // sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                    // sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                   // sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                 // sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                  // sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                 // sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          keys_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                           // keys_s1_translator:uav_waitrequest -> keys_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] keys_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                            // keys_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> keys_s1_translator:uav_burstcount
	wire   [31:0] keys_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                             // keys_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> keys_s1_translator:uav_writedata
	wire   [31:0] keys_s1_translator_avalon_universal_slave_0_agent_m0_address;                                               // keys_s1_translator_avalon_universal_slave_0_agent:m0_address -> keys_s1_translator:uav_address
	wire          keys_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                 // keys_s1_translator_avalon_universal_slave_0_agent:m0_write -> keys_s1_translator:uav_write
	wire          keys_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                  // keys_s1_translator_avalon_universal_slave_0_agent:m0_lock -> keys_s1_translator:uav_lock
	wire          keys_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                  // keys_s1_translator_avalon_universal_slave_0_agent:m0_read -> keys_s1_translator:uav_read
	wire   [31:0] keys_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                              // keys_s1_translator:uav_readdata -> keys_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          keys_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                         // keys_s1_translator:uav_readdatavalid -> keys_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          keys_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                           // keys_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> keys_s1_translator:uav_debugaccess
	wire    [3:0] keys_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                            // keys_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> keys_s1_translator:uav_byteenable
	wire          keys_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                    // keys_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          keys_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                          // keys_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          keys_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                  // keys_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] keys_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                           // keys_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          keys_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                          // keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> keys_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                 // keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> keys_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                       // keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> keys_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                               // keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> keys_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                        // keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> keys_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                       // keys_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          keys_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                     // keys_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> keys_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] keys_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                      // keys_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> keys_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          keys_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                     // keys_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> keys_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          leds_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                           // LEDs_s1_translator:uav_waitrequest -> LEDs_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] leds_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                            // LEDs_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> LEDs_s1_translator:uav_burstcount
	wire   [31:0] leds_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                             // LEDs_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> LEDs_s1_translator:uav_writedata
	wire   [31:0] leds_s1_translator_avalon_universal_slave_0_agent_m0_address;                                               // LEDs_s1_translator_avalon_universal_slave_0_agent:m0_address -> LEDs_s1_translator:uav_address
	wire          leds_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                 // LEDs_s1_translator_avalon_universal_slave_0_agent:m0_write -> LEDs_s1_translator:uav_write
	wire          leds_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                  // LEDs_s1_translator_avalon_universal_slave_0_agent:m0_lock -> LEDs_s1_translator:uav_lock
	wire          leds_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                  // LEDs_s1_translator_avalon_universal_slave_0_agent:m0_read -> LEDs_s1_translator:uav_read
	wire   [31:0] leds_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                              // LEDs_s1_translator:uav_readdata -> LEDs_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          leds_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                         // LEDs_s1_translator:uav_readdatavalid -> LEDs_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          leds_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                           // LEDs_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> LEDs_s1_translator:uav_debugaccess
	wire    [3:0] leds_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                            // LEDs_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> LEDs_s1_translator:uav_byteenable
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                    // LEDs_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> LEDs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                          // LEDs_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> LEDs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                  // LEDs_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> LEDs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] leds_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                           // LEDs_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> LEDs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                          // LEDs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> LEDs_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                 // LEDs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> LEDs_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                       // LEDs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> LEDs_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                               // LEDs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> LEDs_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                        // LEDs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> LEDs_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                       // LEDs_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> LEDs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                     // LEDs_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> LEDs_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                      // LEDs_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> LEDs_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                     // LEDs_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> LEDs_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                     // jtag_uart_0_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                      // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_0_avalon_jtag_slave_translator:uav_burstcount
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                       // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_0_avalon_jtag_slave_translator:uav_writedata
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                         // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_0_avalon_jtag_slave_translator:uav_address
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                           // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_0_avalon_jtag_slave_translator:uav_write
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                            // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_0_avalon_jtag_slave_translator:uav_lock
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                            // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_0_avalon_jtag_slave_translator:uav_read
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                        // jtag_uart_0_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                   // jtag_uart_0_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                     // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_0_avalon_jtag_slave_translator:uav_debugaccess
	wire    [3:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                      // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_0_avalon_jtag_slave_translator:uav_byteenable
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;              // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;            // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                     // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;           // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                 // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;         // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                  // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                 // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;               // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;               // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                  // character_lcd_0_avalon_lcd_slave_translator:uav_waitrequest -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [0:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                   // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> character_lcd_0_avalon_lcd_slave_translator:uav_burstcount
	wire    [7:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                    // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> character_lcd_0_avalon_lcd_slave_translator:uav_writedata
	wire   [31:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_address;                      // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_address -> character_lcd_0_avalon_lcd_slave_translator:uav_address
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_write;                        // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_write -> character_lcd_0_avalon_lcd_slave_translator:uav_write
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_lock;                         // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_lock -> character_lcd_0_avalon_lcd_slave_translator:uav_lock
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_read;                         // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_read -> character_lcd_0_avalon_lcd_slave_translator:uav_read
	wire    [7:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                     // character_lcd_0_avalon_lcd_slave_translator:uav_readdata -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                // character_lcd_0_avalon_lcd_slave_translator:uav_readdatavalid -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                  // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> character_lcd_0_avalon_lcd_slave_translator:uav_debugaccess
	wire    [0:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                   // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> character_lcd_0_avalon_lcd_slave_translator:uav_byteenable
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;           // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                 // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;         // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [80:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                  // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                 // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;        // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;              // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;      // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [80:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;               // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;              // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;            // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire    [9:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;             // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;            // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                    // pixel_buffer_avalon_sram_slave_translator:uav_waitrequest -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [1:0] pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                     // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> pixel_buffer_avalon_sram_slave_translator:uav_burstcount
	wire   [15:0] pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                      // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> pixel_buffer_avalon_sram_slave_translator:uav_writedata
	wire   [31:0] pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address;                        // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_address -> pixel_buffer_avalon_sram_slave_translator:uav_address
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write;                          // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_write -> pixel_buffer_avalon_sram_slave_translator:uav_write
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock;                           // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_lock -> pixel_buffer_avalon_sram_slave_translator:uav_lock
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read;                           // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_read -> pixel_buffer_avalon_sram_slave_translator:uav_read
	wire   [15:0] pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                       // pixel_buffer_avalon_sram_slave_translator:uav_readdata -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                  // pixel_buffer_avalon_sram_slave_translator:uav_readdatavalid -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                    // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pixel_buffer_avalon_sram_slave_translator:uav_debugaccess
	wire    [1:0] pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                     // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> pixel_buffer_avalon_sram_slave_translator:uav_byteenable
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;             // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                   // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;           // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [89:0] pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                    // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                   // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;          // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;        // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [89:0] pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                 // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;              // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [17:0] pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;               // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;              // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;              // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [17:0] pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;               // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;              // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // pixel_buffer_dma_avalon_control_slave_translator:uav_waitrequest -> pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> pixel_buffer_dma_avalon_control_slave_translator:uav_burstcount
	wire   [31:0] pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> pixel_buffer_dma_avalon_control_slave_translator:uav_writedata
	wire   [31:0] pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> pixel_buffer_dma_avalon_control_slave_translator:uav_address
	wire          pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> pixel_buffer_dma_avalon_control_slave_translator:uav_write
	wire          pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> pixel_buffer_dma_avalon_control_slave_translator:uav_lock
	wire          pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> pixel_buffer_dma_avalon_control_slave_translator:uav_read
	wire   [31:0] pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // pixel_buffer_dma_avalon_control_slave_translator:uav_readdata -> pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // pixel_buffer_dma_avalon_control_slave_translator:uav_readdatavalid -> pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pixel_buffer_dma_avalon_control_slave_translator:uav_debugaccess
	wire    [3:0] pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> pixel_buffer_dma_avalon_control_slave_translator:uav_byteenable
	wire          pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                      // line_drawer_0_avalon_slave_0_translator:uav_waitrequest -> line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;                       // line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> line_drawer_0_avalon_slave_0_translator:uav_burstcount
	wire   [31:0] line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;                        // line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> line_drawer_0_avalon_slave_0_translator:uav_writedata
	wire   [31:0] line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                          // line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> line_drawer_0_avalon_slave_0_translator:uav_address
	wire          line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                            // line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> line_drawer_0_avalon_slave_0_translator:uav_write
	wire          line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                             // line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> line_drawer_0_avalon_slave_0_translator:uav_lock
	wire          line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                             // line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> line_drawer_0_avalon_slave_0_translator:uav_read
	wire   [31:0] line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                         // line_drawer_0_avalon_slave_0_translator:uav_readdata -> line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                    // line_drawer_0_avalon_slave_0_translator:uav_readdatavalid -> line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                      // line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> line_drawer_0_avalon_slave_0_translator:uav_debugaccess
	wire    [3:0] line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;                       // line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> line_drawer_0_avalon_slave_0_translator:uav_byteenable
	wire          line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;               // line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;                     // line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;             // line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;                      // line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;                     // line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;            // line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                  // line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;          // line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                   // line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                  // line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                // line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                 // line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                // line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          dual_port_ram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // dual_port_ram_s1_translator:uav_waitrequest -> dual_port_ram_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [0:0] dual_port_ram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // dual_port_ram_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> dual_port_ram_s1_translator:uav_burstcount
	wire    [7:0] dual_port_ram_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // dual_port_ram_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> dual_port_ram_s1_translator:uav_writedata
	wire   [31:0] dual_port_ram_s1_translator_avalon_universal_slave_0_agent_m0_address;                                      // dual_port_ram_s1_translator_avalon_universal_slave_0_agent:m0_address -> dual_port_ram_s1_translator:uav_address
	wire          dual_port_ram_s1_translator_avalon_universal_slave_0_agent_m0_write;                                        // dual_port_ram_s1_translator_avalon_universal_slave_0_agent:m0_write -> dual_port_ram_s1_translator:uav_write
	wire          dual_port_ram_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                         // dual_port_ram_s1_translator_avalon_universal_slave_0_agent:m0_lock -> dual_port_ram_s1_translator:uav_lock
	wire          dual_port_ram_s1_translator_avalon_universal_slave_0_agent_m0_read;                                         // dual_port_ram_s1_translator_avalon_universal_slave_0_agent:m0_read -> dual_port_ram_s1_translator:uav_read
	wire    [7:0] dual_port_ram_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // dual_port_ram_s1_translator:uav_readdata -> dual_port_ram_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          dual_port_ram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // dual_port_ram_s1_translator:uav_readdatavalid -> dual_port_ram_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          dual_port_ram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // dual_port_ram_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> dual_port_ram_s1_translator:uav_debugaccess
	wire    [0:0] dual_port_ram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // dual_port_ram_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> dual_port_ram_s1_translator:uav_byteenable
	wire          dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // dual_port_ram_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // dual_port_ram_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // dual_port_ram_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [80:0] dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // dual_port_ram_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> dual_port_ram_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> dual_port_ram_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> dual_port_ram_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> dual_port_ram_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [80:0] dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> dual_port_ram_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // dual_port_ram_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // dual_port_ram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> dual_port_ram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire    [9:0] dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // dual_port_ram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> dual_port_ram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // dual_port_ram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> dual_port_ram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pi_request_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                     // pi_request_s1_translator:uav_waitrequest -> pi_request_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] pi_request_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                      // pi_request_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pi_request_s1_translator:uav_burstcount
	wire   [31:0] pi_request_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                       // pi_request_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pi_request_s1_translator:uav_writedata
	wire   [31:0] pi_request_s1_translator_avalon_universal_slave_0_agent_m0_address;                                         // pi_request_s1_translator_avalon_universal_slave_0_agent:m0_address -> pi_request_s1_translator:uav_address
	wire          pi_request_s1_translator_avalon_universal_slave_0_agent_m0_write;                                           // pi_request_s1_translator_avalon_universal_slave_0_agent:m0_write -> pi_request_s1_translator:uav_write
	wire          pi_request_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                            // pi_request_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pi_request_s1_translator:uav_lock
	wire          pi_request_s1_translator_avalon_universal_slave_0_agent_m0_read;                                            // pi_request_s1_translator_avalon_universal_slave_0_agent:m0_read -> pi_request_s1_translator:uav_read
	wire   [31:0] pi_request_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                        // pi_request_s1_translator:uav_readdata -> pi_request_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          pi_request_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                   // pi_request_s1_translator:uav_readdatavalid -> pi_request_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          pi_request_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                     // pi_request_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pi_request_s1_translator:uav_debugaccess
	wire    [3:0] pi_request_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                      // pi_request_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pi_request_s1_translator:uav_byteenable
	wire          pi_request_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                              // pi_request_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pi_request_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          pi_request_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                    // pi_request_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pi_request_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          pi_request_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                            // pi_request_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pi_request_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] pi_request_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                     // pi_request_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pi_request_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          pi_request_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                    // pi_request_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pi_request_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          pi_request_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                           // pi_request_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pi_request_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          pi_request_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                 // pi_request_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pi_request_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          pi_request_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                         // pi_request_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pi_request_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] pi_request_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                  // pi_request_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pi_request_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          pi_request_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                 // pi_request_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pi_request_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          pi_request_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                               // pi_request_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pi_request_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] pi_request_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                // pi_request_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pi_request_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          pi_request_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                               // pi_request_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pi_request_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          de2_ack_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                        // de2_ack_s1_translator:uav_waitrequest -> de2_ack_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] de2_ack_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                         // de2_ack_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> de2_ack_s1_translator:uav_burstcount
	wire   [31:0] de2_ack_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                          // de2_ack_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> de2_ack_s1_translator:uav_writedata
	wire   [31:0] de2_ack_s1_translator_avalon_universal_slave_0_agent_m0_address;                                            // de2_ack_s1_translator_avalon_universal_slave_0_agent:m0_address -> de2_ack_s1_translator:uav_address
	wire          de2_ack_s1_translator_avalon_universal_slave_0_agent_m0_write;                                              // de2_ack_s1_translator_avalon_universal_slave_0_agent:m0_write -> de2_ack_s1_translator:uav_write
	wire          de2_ack_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                               // de2_ack_s1_translator_avalon_universal_slave_0_agent:m0_lock -> de2_ack_s1_translator:uav_lock
	wire          de2_ack_s1_translator_avalon_universal_slave_0_agent_m0_read;                                               // de2_ack_s1_translator_avalon_universal_slave_0_agent:m0_read -> de2_ack_s1_translator:uav_read
	wire   [31:0] de2_ack_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                           // de2_ack_s1_translator:uav_readdata -> de2_ack_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          de2_ack_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                      // de2_ack_s1_translator:uav_readdatavalid -> de2_ack_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          de2_ack_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                        // de2_ack_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> de2_ack_s1_translator:uav_debugaccess
	wire    [3:0] de2_ack_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                         // de2_ack_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> de2_ack_s1_translator:uav_byteenable
	wire          de2_ack_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                 // de2_ack_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> de2_ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          de2_ack_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                       // de2_ack_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> de2_ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          de2_ack_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                               // de2_ack_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> de2_ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] de2_ack_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                        // de2_ack_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> de2_ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          de2_ack_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                       // de2_ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> de2_ack_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          de2_ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                              // de2_ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> de2_ack_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          de2_ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                    // de2_ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> de2_ack_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          de2_ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                            // de2_ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> de2_ack_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] de2_ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                     // de2_ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> de2_ack_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          de2_ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                    // de2_ack_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> de2_ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          de2_ack_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                  // de2_ack_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> de2_ack_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] de2_ack_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                   // de2_ack_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> de2_ack_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          de2_ack_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                  // de2_ack_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> de2_ack_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                  // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire          nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                        // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire          nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [106:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                         // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire          nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                        // addr_router:sink_ready -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                         // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire          nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_valid;                               // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire          nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                       // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [106:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_data;                                // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire          nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_ready;                               // addr_router_001:sink_ready -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket;         // pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_002:sink_endofpacket
	wire          pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_valid;               // pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_002:sink_valid
	wire          pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket;       // pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_002:sink_startofpacket
	wire   [88:0] pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_data;                // pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_002:sink_data
	wire          pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_ready;               // addr_router_002:sink_ready -> pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          line_drawer_0_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                      // line_drawer_0_avalon_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_003:sink_endofpacket
	wire          line_drawer_0_avalon_master_translator_avalon_universal_master_0_agent_cp_valid;                            // line_drawer_0_avalon_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_003:sink_valid
	wire          line_drawer_0_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                    // line_drawer_0_avalon_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_003:sink_startofpacket
	wire   [88:0] line_drawer_0_avalon_master_translator_avalon_universal_master_0_agent_cp_data;                             // line_drawer_0_avalon_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_003:sink_data
	wire          line_drawer_0_avalon_master_translator_avalon_universal_master_0_agent_cp_ready;                            // addr_router_003:sink_ready -> line_drawer_0_avalon_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                    // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                          // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                  // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [106:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                           // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                          // id_router:sink_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                     // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [106:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                      // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_001:sink_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                          // sdram_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                // sdram_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                        // sdram_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire   [88:0] sdram_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                 // sdram_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                // id_router_002:sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          timer_system_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                   // timer_system_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire          timer_system_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                         // timer_system_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire          timer_system_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                 // timer_system_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [106:0] timer_system_s1_translator_avalon_universal_slave_0_agent_rp_data;                                          // timer_system_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire          timer_system_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                         // id_router_003:sink_ready -> timer_system_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // timer_timestamp_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire          timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                      // timer_timestamp_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire          timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // timer_timestamp_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [106:0] timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rp_data;                                       // timer_timestamp_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire          timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_004:sink_ready -> timer_timestamp_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                       // sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_valid;                             // sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                     // sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [106:0] sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_data;                              // sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_ready;                             // id_router_005:sink_ready -> sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          keys_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                           // keys_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire          keys_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                 // keys_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire          keys_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                         // keys_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire  [106:0] keys_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                  // keys_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire          keys_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                 // id_router_006:sink_ready -> keys_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                           // LEDs_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                 // LEDs_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                         // LEDs_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire  [106:0] leds_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                  // LEDs_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                 // id_router_007:sink_ready -> LEDs_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                     // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                           // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                   // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire  [106:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                            // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                           // id_router_008:sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                  // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_valid;                        // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	wire   [79:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_data;                         // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_ready;                        // id_router_009:sink_ready -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                    // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid;                          // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                  // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	wire   [88:0] pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data;                           // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready;                          // id_router_010:sink_ready -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	wire          pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	wire          pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	wire  [106:0] pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	wire          pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_011:sink_ready -> pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                      // line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	wire          line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                            // line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	wire          line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                    // line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	wire  [106:0] line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                             // line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	wire          line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                            // id_router_012:sink_ready -> line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // dual_port_ram_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_013:sink_endofpacket
	wire          dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                        // dual_port_ram_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_013:sink_valid
	wire          dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // dual_port_ram_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_013:sink_startofpacket
	wire   [79:0] dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rp_data;                                         // dual_port_ram_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_013:sink_data
	wire          dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_013:sink_ready -> dual_port_ram_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pi_request_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                     // pi_request_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_014:sink_endofpacket
	wire          pi_request_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                           // pi_request_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_014:sink_valid
	wire          pi_request_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                   // pi_request_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_014:sink_startofpacket
	wire  [106:0] pi_request_s1_translator_avalon_universal_slave_0_agent_rp_data;                                            // pi_request_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_014:sink_data
	wire          pi_request_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                           // id_router_014:sink_ready -> pi_request_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          de2_ack_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                        // de2_ack_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_015:sink_endofpacket
	wire          de2_ack_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                              // de2_ack_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_015:sink_valid
	wire          de2_ack_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                      // de2_ack_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_015:sink_startofpacket
	wire  [106:0] de2_ack_s1_translator_avalon_universal_slave_0_agent_rp_data;                                               // de2_ack_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_015:sink_data
	wire          de2_ack_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                              // id_router_015:sink_ready -> de2_ack_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          burst_adapter_source0_endofpacket;                                                                          // burst_adapter:source0_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_source0_valid;                                                                                // burst_adapter:source0_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_source0_startofpacket;                                                                        // burst_adapter:source0_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [88:0] burst_adapter_source0_data;                                                                                 // burst_adapter:source0_data -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_source0_ready;                                                                                // sdram_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	wire   [15:0] burst_adapter_source0_channel;                                                                              // burst_adapter:source0_channel -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_001_source0_endofpacket;                                                                      // burst_adapter_001:source0_endofpacket -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_001_source0_valid;                                                                            // burst_adapter_001:source0_valid -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_001_source0_startofpacket;                                                                    // burst_adapter_001:source0_startofpacket -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [79:0] burst_adapter_001_source0_data;                                                                             // burst_adapter_001:source0_data -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_001_source0_ready;                                                                            // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_001:source0_ready
	wire   [15:0] burst_adapter_001_source0_channel;                                                                          // burst_adapter_001:source0_channel -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_002_source0_endofpacket;                                                                      // burst_adapter_002:source0_endofpacket -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_002_source0_valid;                                                                            // burst_adapter_002:source0_valid -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_002_source0_startofpacket;                                                                    // burst_adapter_002:source0_startofpacket -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [88:0] burst_adapter_002_source0_data;                                                                             // burst_adapter_002:source0_data -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_002_source0_ready;                                                                            // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_002:source0_ready
	wire   [15:0] burst_adapter_002_source0_channel;                                                                          // burst_adapter_002:source0_channel -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_003_source0_endofpacket;                                                                      // burst_adapter_003:source0_endofpacket -> dual_port_ram_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_003_source0_valid;                                                                            // burst_adapter_003:source0_valid -> dual_port_ram_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_003_source0_startofpacket;                                                                    // burst_adapter_003:source0_startofpacket -> dual_port_ram_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [79:0] burst_adapter_003_source0_data;                                                                             // burst_adapter_003:source0_data -> dual_port_ram_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_003_source0_ready;                                                                            // dual_port_ram_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_003:source0_ready
	wire   [15:0] burst_adapter_003_source0_channel;                                                                          // burst_adapter_003:source0_channel -> dual_port_ram_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rst_controller_reset_out_reset;                                                                             // rst_controller:reset_out -> [LEDs:reset_n, LEDs_s1_translator:reset, LEDs_s1_translator_avalon_universal_slave_0_agent:reset, LEDs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, addr_router:reset, addr_router_001:reset, addr_router_002:reset, addr_router_003:reset, burst_adapter:reset, burst_adapter_001:reset, burst_adapter_002:reset, burst_adapter_003:reset, character_lcd_0:reset, character_lcd_0_avalon_lcd_slave_translator:reset, character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:reset, character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_demux_002:reset, cmd_xbar_demux_003:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_002:reset, cmd_xbar_mux_003:reset, cmd_xbar_mux_004:reset, cmd_xbar_mux_005:reset, cmd_xbar_mux_010:reset, de2_ack:reset_n, de2_ack_s1_translator:reset, de2_ack_s1_translator_avalon_universal_slave_0_agent:reset, de2_ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, dual_port_ram:reset, dual_port_ram_s1_translator:reset, dual_port_ram_s1_translator_avalon_universal_slave_0_agent:reset, dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_010:reset, id_router_011:reset, id_router_012:reset, id_router_013:reset, id_router_014:reset, id_router_015:reset, irq_mapper:reset, jtag_uart_0:rst_n, jtag_uart_0_avalon_jtag_slave_translator:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, keys:reset_n, keys_s1_translator:reset, keys_s1_translator_avalon_universal_slave_0_agent:reset, keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, line_drawer_0:reset_n, line_drawer_0_avalon_master_translator:reset, line_drawer_0_avalon_master_translator_avalon_universal_master_0_agent:reset, line_drawer_0_avalon_slave_0_translator:reset, line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, nios2_qsys_0:reset_n, nios2_qsys_0_data_master_translator:reset, nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:reset, nios2_qsys_0_instruction_master_translator:reset, nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:reset, nios2_qsys_0_jtag_debug_module_translator:reset, nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, onchip_memory2_0:reset, onchip_memory2_0_s1_translator:reset, onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:reset, onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pi_request:reset_n, pi_request_s1_translator:reset, pi_request_s1_translator_avalon_universal_slave_0_agent:reset, pi_request_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pixel_buffer:reset, pixel_buffer_avalon_sram_slave_translator:reset, pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:reset, pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pixel_buffer_dma:reset, pixel_buffer_dma_avalon_control_slave_translator:reset, pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:reset, pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pixel_buffer_dma_avalon_pixel_dma_master_translator:reset, pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:reset, rgb_sampler:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset, rsp_xbar_demux_011:reset, rsp_xbar_demux_012:reset, rsp_xbar_demux_013:reset, rsp_xbar_demux_014:reset, rsp_xbar_demux_015:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, scaler:reset, sd_card:i_reset_n, sd_card_avalon_sdcard_slave_translator:reset, sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:reset, sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sdram:reset_n, sdram_s1_translator:reset, sdram_s1_translator_avalon_universal_slave_0_agent:reset, sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timer_system:reset_n, timer_system_s1_translator:reset, timer_system_s1_translator_avalon_universal_slave_0_agent:reset, timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timer_timestamp:reset_n, timer_timestamp_s1_translator:reset, timer_timestamp_s1_translator_avalon_universal_slave_0_agent:reset, timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, video_fifo:reset_stream_in, width_adapter:reset, width_adapter_001:reset, width_adapter_002:reset, width_adapter_003:reset, width_adapter_004:reset, width_adapter_005:reset, width_adapter_006:reset, width_adapter_007:reset, width_adapter_008:reset, width_adapter_009:reset]
	wire          rst_controller_reset_out_reset_req;                                                                         // rst_controller:reset_req -> [dual_port_ram:reset_req, onchip_memory2_0:reset_req]
	wire          nios2_qsys_0_jtag_debug_module_reset_reset;                                                                 // nios2_qsys_0:jtag_debug_module_resetrequest -> [rst_controller:reset_in0, rst_controller_001:reset_in1, rst_controller_002:reset_in1, rst_controller_003:reset_in1, rst_controller_004:reset_in0]
	wire          rst_controller_001_reset_out_reset;                                                                         // rst_controller_001:reset_out -> clocks:reset
	wire          rst_controller_002_reset_out_reset;                                                                         // rst_controller_002:reset_out -> [vga_controller:reset, video_fifo:reset_stream_out]
	wire          rst_controller_003_reset_out_reset;                                                                         // rst_controller_003:reset_out -> dual_port_ram:reset2
	wire          rst_controller_003_reset_out_reset_req;                                                                     // rst_controller_003:reset_req -> dual_port_ram:reset_req2
	wire          rst_controller_004_reset_out_reset;                                                                         // rst_controller_004:reset_out -> rst_controller_003:reset_in2
	wire          cmd_xbar_demux_src0_endofpacket;                                                                            // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                                                                  // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                                                          // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_src0_data;                                                                                   // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire   [15:0] cmd_xbar_demux_src0_channel;                                                                                // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire          cmd_xbar_demux_src0_ready;                                                                                  // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire          cmd_xbar_demux_src1_endofpacket;                                                                            // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire          cmd_xbar_demux_src1_valid;                                                                                  // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire          cmd_xbar_demux_src1_startofpacket;                                                                          // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_src1_data;                                                                                   // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire   [15:0] cmd_xbar_demux_src1_channel;                                                                                // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire          cmd_xbar_demux_src1_ready;                                                                                  // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire          cmd_xbar_demux_src3_endofpacket;                                                                            // cmd_xbar_demux:src3_endofpacket -> cmd_xbar_mux_003:sink0_endofpacket
	wire          cmd_xbar_demux_src3_valid;                                                                                  // cmd_xbar_demux:src3_valid -> cmd_xbar_mux_003:sink0_valid
	wire          cmd_xbar_demux_src3_startofpacket;                                                                          // cmd_xbar_demux:src3_startofpacket -> cmd_xbar_mux_003:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_src3_data;                                                                                   // cmd_xbar_demux:src3_data -> cmd_xbar_mux_003:sink0_data
	wire   [15:0] cmd_xbar_demux_src3_channel;                                                                                // cmd_xbar_demux:src3_channel -> cmd_xbar_mux_003:sink0_channel
	wire          cmd_xbar_demux_src3_ready;                                                                                  // cmd_xbar_mux_003:sink0_ready -> cmd_xbar_demux:src3_ready
	wire          cmd_xbar_demux_src4_endofpacket;                                                                            // cmd_xbar_demux:src4_endofpacket -> cmd_xbar_mux_004:sink0_endofpacket
	wire          cmd_xbar_demux_src4_valid;                                                                                  // cmd_xbar_demux:src4_valid -> cmd_xbar_mux_004:sink0_valid
	wire          cmd_xbar_demux_src4_startofpacket;                                                                          // cmd_xbar_demux:src4_startofpacket -> cmd_xbar_mux_004:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_src4_data;                                                                                   // cmd_xbar_demux:src4_data -> cmd_xbar_mux_004:sink0_data
	wire   [15:0] cmd_xbar_demux_src4_channel;                                                                                // cmd_xbar_demux:src4_channel -> cmd_xbar_mux_004:sink0_channel
	wire          cmd_xbar_demux_src4_ready;                                                                                  // cmd_xbar_mux_004:sink0_ready -> cmd_xbar_demux:src4_ready
	wire          cmd_xbar_demux_src5_endofpacket;                                                                            // cmd_xbar_demux:src5_endofpacket -> cmd_xbar_mux_005:sink0_endofpacket
	wire          cmd_xbar_demux_src5_valid;                                                                                  // cmd_xbar_demux:src5_valid -> cmd_xbar_mux_005:sink0_valid
	wire          cmd_xbar_demux_src5_startofpacket;                                                                          // cmd_xbar_demux:src5_startofpacket -> cmd_xbar_mux_005:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_src5_data;                                                                                   // cmd_xbar_demux:src5_data -> cmd_xbar_mux_005:sink0_data
	wire   [15:0] cmd_xbar_demux_src5_channel;                                                                                // cmd_xbar_demux:src5_channel -> cmd_xbar_mux_005:sink0_channel
	wire          cmd_xbar_demux_src5_ready;                                                                                  // cmd_xbar_mux_005:sink0_ready -> cmd_xbar_demux:src5_ready
	wire          cmd_xbar_demux_001_src0_endofpacket;                                                                        // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire          cmd_xbar_demux_001_src0_valid;                                                                              // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire          cmd_xbar_demux_001_src0_startofpacket;                                                                      // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src0_data;                                                                               // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire   [15:0] cmd_xbar_demux_001_src0_channel;                                                                            // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire          cmd_xbar_demux_001_src0_ready;                                                                              // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire          cmd_xbar_demux_001_src1_endofpacket;                                                                        // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire          cmd_xbar_demux_001_src1_valid;                                                                              // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	wire          cmd_xbar_demux_001_src1_startofpacket;                                                                      // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src1_data;                                                                               // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	wire   [15:0] cmd_xbar_demux_001_src1_channel;                                                                            // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	wire          cmd_xbar_demux_001_src1_ready;                                                                              // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire          cmd_xbar_demux_001_src3_endofpacket;                                                                        // cmd_xbar_demux_001:src3_endofpacket -> cmd_xbar_mux_003:sink1_endofpacket
	wire          cmd_xbar_demux_001_src3_valid;                                                                              // cmd_xbar_demux_001:src3_valid -> cmd_xbar_mux_003:sink1_valid
	wire          cmd_xbar_demux_001_src3_startofpacket;                                                                      // cmd_xbar_demux_001:src3_startofpacket -> cmd_xbar_mux_003:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src3_data;                                                                               // cmd_xbar_demux_001:src3_data -> cmd_xbar_mux_003:sink1_data
	wire   [15:0] cmd_xbar_demux_001_src3_channel;                                                                            // cmd_xbar_demux_001:src3_channel -> cmd_xbar_mux_003:sink1_channel
	wire          cmd_xbar_demux_001_src3_ready;                                                                              // cmd_xbar_mux_003:sink1_ready -> cmd_xbar_demux_001:src3_ready
	wire          cmd_xbar_demux_001_src4_endofpacket;                                                                        // cmd_xbar_demux_001:src4_endofpacket -> cmd_xbar_mux_004:sink1_endofpacket
	wire          cmd_xbar_demux_001_src4_valid;                                                                              // cmd_xbar_demux_001:src4_valid -> cmd_xbar_mux_004:sink1_valid
	wire          cmd_xbar_demux_001_src4_startofpacket;                                                                      // cmd_xbar_demux_001:src4_startofpacket -> cmd_xbar_mux_004:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src4_data;                                                                               // cmd_xbar_demux_001:src4_data -> cmd_xbar_mux_004:sink1_data
	wire   [15:0] cmd_xbar_demux_001_src4_channel;                                                                            // cmd_xbar_demux_001:src4_channel -> cmd_xbar_mux_004:sink1_channel
	wire          cmd_xbar_demux_001_src4_ready;                                                                              // cmd_xbar_mux_004:sink1_ready -> cmd_xbar_demux_001:src4_ready
	wire          cmd_xbar_demux_001_src5_endofpacket;                                                                        // cmd_xbar_demux_001:src5_endofpacket -> cmd_xbar_mux_005:sink1_endofpacket
	wire          cmd_xbar_demux_001_src5_valid;                                                                              // cmd_xbar_demux_001:src5_valid -> cmd_xbar_mux_005:sink1_valid
	wire          cmd_xbar_demux_001_src5_startofpacket;                                                                      // cmd_xbar_demux_001:src5_startofpacket -> cmd_xbar_mux_005:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src5_data;                                                                               // cmd_xbar_demux_001:src5_data -> cmd_xbar_mux_005:sink1_data
	wire   [15:0] cmd_xbar_demux_001_src5_channel;                                                                            // cmd_xbar_demux_001:src5_channel -> cmd_xbar_mux_005:sink1_channel
	wire          cmd_xbar_demux_001_src5_ready;                                                                              // cmd_xbar_mux_005:sink1_ready -> cmd_xbar_demux_001:src5_ready
	wire          cmd_xbar_demux_001_src6_endofpacket;                                                                        // cmd_xbar_demux_001:src6_endofpacket -> keys_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src6_valid;                                                                              // cmd_xbar_demux_001:src6_valid -> keys_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src6_startofpacket;                                                                      // cmd_xbar_demux_001:src6_startofpacket -> keys_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src6_data;                                                                               // cmd_xbar_demux_001:src6_data -> keys_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_001_src6_channel;                                                                            // cmd_xbar_demux_001:src6_channel -> keys_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src7_endofpacket;                                                                        // cmd_xbar_demux_001:src7_endofpacket -> LEDs_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src7_valid;                                                                              // cmd_xbar_demux_001:src7_valid -> LEDs_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src7_startofpacket;                                                                      // cmd_xbar_demux_001:src7_startofpacket -> LEDs_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src7_data;                                                                               // cmd_xbar_demux_001:src7_data -> LEDs_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_001_src7_channel;                                                                            // cmd_xbar_demux_001:src7_channel -> LEDs_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src8_endofpacket;                                                                        // cmd_xbar_demux_001:src8_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src8_valid;                                                                              // cmd_xbar_demux_001:src8_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src8_startofpacket;                                                                      // cmd_xbar_demux_001:src8_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src8_data;                                                                               // cmd_xbar_demux_001:src8_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_001_src8_channel;                                                                            // cmd_xbar_demux_001:src8_channel -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src11_endofpacket;                                                                       // cmd_xbar_demux_001:src11_endofpacket -> pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src11_valid;                                                                             // cmd_xbar_demux_001:src11_valid -> pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src11_startofpacket;                                                                     // cmd_xbar_demux_001:src11_startofpacket -> pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src11_data;                                                                              // cmd_xbar_demux_001:src11_data -> pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_001_src11_channel;                                                                           // cmd_xbar_demux_001:src11_channel -> pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src12_endofpacket;                                                                       // cmd_xbar_demux_001:src12_endofpacket -> line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src12_valid;                                                                             // cmd_xbar_demux_001:src12_valid -> line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src12_startofpacket;                                                                     // cmd_xbar_demux_001:src12_startofpacket -> line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src12_data;                                                                              // cmd_xbar_demux_001:src12_data -> line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_001_src12_channel;                                                                           // cmd_xbar_demux_001:src12_channel -> line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src14_endofpacket;                                                                       // cmd_xbar_demux_001:src14_endofpacket -> pi_request_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src14_valid;                                                                             // cmd_xbar_demux_001:src14_valid -> pi_request_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src14_startofpacket;                                                                     // cmd_xbar_demux_001:src14_startofpacket -> pi_request_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src14_data;                                                                              // cmd_xbar_demux_001:src14_data -> pi_request_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_001_src14_channel;                                                                           // cmd_xbar_demux_001:src14_channel -> pi_request_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src15_endofpacket;                                                                       // cmd_xbar_demux_001:src15_endofpacket -> de2_ack_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src15_valid;                                                                             // cmd_xbar_demux_001:src15_valid -> de2_ack_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src15_startofpacket;                                                                     // cmd_xbar_demux_001:src15_startofpacket -> de2_ack_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src15_data;                                                                              // cmd_xbar_demux_001:src15_data -> de2_ack_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_001_src15_channel;                                                                           // cmd_xbar_demux_001:src15_channel -> de2_ack_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_002_src0_endofpacket;                                                                        // cmd_xbar_demux_002:src0_endofpacket -> cmd_xbar_mux_010:sink1_endofpacket
	wire          cmd_xbar_demux_002_src0_valid;                                                                              // cmd_xbar_demux_002:src0_valid -> cmd_xbar_mux_010:sink1_valid
	wire          cmd_xbar_demux_002_src0_startofpacket;                                                                      // cmd_xbar_demux_002:src0_startofpacket -> cmd_xbar_mux_010:sink1_startofpacket
	wire   [88:0] cmd_xbar_demux_002_src0_data;                                                                               // cmd_xbar_demux_002:src0_data -> cmd_xbar_mux_010:sink1_data
	wire   [15:0] cmd_xbar_demux_002_src0_channel;                                                                            // cmd_xbar_demux_002:src0_channel -> cmd_xbar_mux_010:sink1_channel
	wire          cmd_xbar_demux_002_src0_ready;                                                                              // cmd_xbar_mux_010:sink1_ready -> cmd_xbar_demux_002:src0_ready
	wire          cmd_xbar_demux_003_src0_endofpacket;                                                                        // cmd_xbar_demux_003:src0_endofpacket -> cmd_xbar_mux_010:sink2_endofpacket
	wire          cmd_xbar_demux_003_src0_valid;                                                                              // cmd_xbar_demux_003:src0_valid -> cmd_xbar_mux_010:sink2_valid
	wire          cmd_xbar_demux_003_src0_startofpacket;                                                                      // cmd_xbar_demux_003:src0_startofpacket -> cmd_xbar_mux_010:sink2_startofpacket
	wire   [88:0] cmd_xbar_demux_003_src0_data;                                                                               // cmd_xbar_demux_003:src0_data -> cmd_xbar_mux_010:sink2_data
	wire   [15:0] cmd_xbar_demux_003_src0_channel;                                                                            // cmd_xbar_demux_003:src0_channel -> cmd_xbar_mux_010:sink2_channel
	wire          cmd_xbar_demux_003_src0_ready;                                                                              // cmd_xbar_mux_010:sink2_ready -> cmd_xbar_demux_003:src0_ready
	wire          rsp_xbar_demux_src0_endofpacket;                                                                            // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                                                                  // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                                                          // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [106:0] rsp_xbar_demux_src0_data;                                                                                   // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire   [15:0] rsp_xbar_demux_src0_channel;                                                                                // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire          rsp_xbar_demux_src0_ready;                                                                                  // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire          rsp_xbar_demux_src1_endofpacket;                                                                            // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire          rsp_xbar_demux_src1_valid;                                                                                  // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire          rsp_xbar_demux_src1_startofpacket;                                                                          // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [106:0] rsp_xbar_demux_src1_data;                                                                                   // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire   [15:0] rsp_xbar_demux_src1_channel;                                                                                // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire          rsp_xbar_demux_src1_ready;                                                                                  // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire          rsp_xbar_demux_001_src0_endofpacket;                                                                        // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire          rsp_xbar_demux_001_src0_valid;                                                                              // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire          rsp_xbar_demux_001_src0_startofpacket;                                                                      // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [106:0] rsp_xbar_demux_001_src0_data;                                                                               // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire   [15:0] rsp_xbar_demux_001_src0_channel;                                                                            // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire          rsp_xbar_demux_001_src0_ready;                                                                              // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire          rsp_xbar_demux_001_src1_endofpacket;                                                                        // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire          rsp_xbar_demux_001_src1_valid;                                                                              // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire          rsp_xbar_demux_001_src1_startofpacket;                                                                      // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [106:0] rsp_xbar_demux_001_src1_data;                                                                               // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	wire   [15:0] rsp_xbar_demux_001_src1_channel;                                                                            // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire          rsp_xbar_demux_001_src1_ready;                                                                              // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	wire          rsp_xbar_demux_003_src0_endofpacket;                                                                        // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux:sink3_endofpacket
	wire          rsp_xbar_demux_003_src0_valid;                                                                              // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux:sink3_valid
	wire          rsp_xbar_demux_003_src0_startofpacket;                                                                      // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux:sink3_startofpacket
	wire  [106:0] rsp_xbar_demux_003_src0_data;                                                                               // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux:sink3_data
	wire   [15:0] rsp_xbar_demux_003_src0_channel;                                                                            // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux:sink3_channel
	wire          rsp_xbar_demux_003_src0_ready;                                                                              // rsp_xbar_mux:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire          rsp_xbar_demux_003_src1_endofpacket;                                                                        // rsp_xbar_demux_003:src1_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire          rsp_xbar_demux_003_src1_valid;                                                                              // rsp_xbar_demux_003:src1_valid -> rsp_xbar_mux_001:sink3_valid
	wire          rsp_xbar_demux_003_src1_startofpacket;                                                                      // rsp_xbar_demux_003:src1_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire  [106:0] rsp_xbar_demux_003_src1_data;                                                                               // rsp_xbar_demux_003:src1_data -> rsp_xbar_mux_001:sink3_data
	wire   [15:0] rsp_xbar_demux_003_src1_channel;                                                                            // rsp_xbar_demux_003:src1_channel -> rsp_xbar_mux_001:sink3_channel
	wire          rsp_xbar_demux_003_src1_ready;                                                                              // rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src1_ready
	wire          rsp_xbar_demux_004_src0_endofpacket;                                                                        // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux:sink4_endofpacket
	wire          rsp_xbar_demux_004_src0_valid;                                                                              // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux:sink4_valid
	wire          rsp_xbar_demux_004_src0_startofpacket;                                                                      // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux:sink4_startofpacket
	wire  [106:0] rsp_xbar_demux_004_src0_data;                                                                               // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux:sink4_data
	wire   [15:0] rsp_xbar_demux_004_src0_channel;                                                                            // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux:sink4_channel
	wire          rsp_xbar_demux_004_src0_ready;                                                                              // rsp_xbar_mux:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire          rsp_xbar_demux_004_src1_endofpacket;                                                                        // rsp_xbar_demux_004:src1_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire          rsp_xbar_demux_004_src1_valid;                                                                              // rsp_xbar_demux_004:src1_valid -> rsp_xbar_mux_001:sink4_valid
	wire          rsp_xbar_demux_004_src1_startofpacket;                                                                      // rsp_xbar_demux_004:src1_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire  [106:0] rsp_xbar_demux_004_src1_data;                                                                               // rsp_xbar_demux_004:src1_data -> rsp_xbar_mux_001:sink4_data
	wire   [15:0] rsp_xbar_demux_004_src1_channel;                                                                            // rsp_xbar_demux_004:src1_channel -> rsp_xbar_mux_001:sink4_channel
	wire          rsp_xbar_demux_004_src1_ready;                                                                              // rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src1_ready
	wire          rsp_xbar_demux_005_src0_endofpacket;                                                                        // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux:sink5_endofpacket
	wire          rsp_xbar_demux_005_src0_valid;                                                                              // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux:sink5_valid
	wire          rsp_xbar_demux_005_src0_startofpacket;                                                                      // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux:sink5_startofpacket
	wire  [106:0] rsp_xbar_demux_005_src0_data;                                                                               // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux:sink5_data
	wire   [15:0] rsp_xbar_demux_005_src0_channel;                                                                            // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux:sink5_channel
	wire          rsp_xbar_demux_005_src0_ready;                                                                              // rsp_xbar_mux:sink5_ready -> rsp_xbar_demux_005:src0_ready
	wire          rsp_xbar_demux_005_src1_endofpacket;                                                                        // rsp_xbar_demux_005:src1_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	wire          rsp_xbar_demux_005_src1_valid;                                                                              // rsp_xbar_demux_005:src1_valid -> rsp_xbar_mux_001:sink5_valid
	wire          rsp_xbar_demux_005_src1_startofpacket;                                                                      // rsp_xbar_demux_005:src1_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	wire  [106:0] rsp_xbar_demux_005_src1_data;                                                                               // rsp_xbar_demux_005:src1_data -> rsp_xbar_mux_001:sink5_data
	wire   [15:0] rsp_xbar_demux_005_src1_channel;                                                                            // rsp_xbar_demux_005:src1_channel -> rsp_xbar_mux_001:sink5_channel
	wire          rsp_xbar_demux_005_src1_ready;                                                                              // rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src1_ready
	wire          rsp_xbar_demux_006_src0_endofpacket;                                                                        // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	wire          rsp_xbar_demux_006_src0_valid;                                                                              // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux_001:sink6_valid
	wire          rsp_xbar_demux_006_src0_startofpacket;                                                                      // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	wire  [106:0] rsp_xbar_demux_006_src0_data;                                                                               // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux_001:sink6_data
	wire   [15:0] rsp_xbar_demux_006_src0_channel;                                                                            // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux_001:sink6_channel
	wire          rsp_xbar_demux_006_src0_ready;                                                                              // rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_006:src0_ready
	wire          rsp_xbar_demux_007_src0_endofpacket;                                                                        // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	wire          rsp_xbar_demux_007_src0_valid;                                                                              // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux_001:sink7_valid
	wire          rsp_xbar_demux_007_src0_startofpacket;                                                                      // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	wire  [106:0] rsp_xbar_demux_007_src0_data;                                                                               // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux_001:sink7_data
	wire   [15:0] rsp_xbar_demux_007_src0_channel;                                                                            // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux_001:sink7_channel
	wire          rsp_xbar_demux_007_src0_ready;                                                                              // rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_007:src0_ready
	wire          rsp_xbar_demux_008_src0_endofpacket;                                                                        // rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux_001:sink8_endofpacket
	wire          rsp_xbar_demux_008_src0_valid;                                                                              // rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux_001:sink8_valid
	wire          rsp_xbar_demux_008_src0_startofpacket;                                                                      // rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux_001:sink8_startofpacket
	wire  [106:0] rsp_xbar_demux_008_src0_data;                                                                               // rsp_xbar_demux_008:src0_data -> rsp_xbar_mux_001:sink8_data
	wire   [15:0] rsp_xbar_demux_008_src0_channel;                                                                            // rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux_001:sink8_channel
	wire          rsp_xbar_demux_008_src0_ready;                                                                              // rsp_xbar_mux_001:sink8_ready -> rsp_xbar_demux_008:src0_ready
	wire          rsp_xbar_demux_010_src1_endofpacket;                                                                        // rsp_xbar_demux_010:src1_endofpacket -> pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_010_src1_valid;                                                                              // rsp_xbar_demux_010:src1_valid -> pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_010_src1_startofpacket;                                                                      // rsp_xbar_demux_010:src1_startofpacket -> pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [88:0] rsp_xbar_demux_010_src1_data;                                                                               // rsp_xbar_demux_010:src1_data -> pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [15:0] rsp_xbar_demux_010_src1_channel;                                                                            // rsp_xbar_demux_010:src1_channel -> pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_010_src2_endofpacket;                                                                        // rsp_xbar_demux_010:src2_endofpacket -> line_drawer_0_avalon_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_010_src2_valid;                                                                              // rsp_xbar_demux_010:src2_valid -> line_drawer_0_avalon_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_010_src2_startofpacket;                                                                      // rsp_xbar_demux_010:src2_startofpacket -> line_drawer_0_avalon_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [88:0] rsp_xbar_demux_010_src2_data;                                                                               // rsp_xbar_demux_010:src2_data -> line_drawer_0_avalon_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [15:0] rsp_xbar_demux_010_src2_channel;                                                                            // rsp_xbar_demux_010:src2_channel -> line_drawer_0_avalon_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_011_src0_endofpacket;                                                                        // rsp_xbar_demux_011:src0_endofpacket -> rsp_xbar_mux_001:sink11_endofpacket
	wire          rsp_xbar_demux_011_src0_valid;                                                                              // rsp_xbar_demux_011:src0_valid -> rsp_xbar_mux_001:sink11_valid
	wire          rsp_xbar_demux_011_src0_startofpacket;                                                                      // rsp_xbar_demux_011:src0_startofpacket -> rsp_xbar_mux_001:sink11_startofpacket
	wire  [106:0] rsp_xbar_demux_011_src0_data;                                                                               // rsp_xbar_demux_011:src0_data -> rsp_xbar_mux_001:sink11_data
	wire   [15:0] rsp_xbar_demux_011_src0_channel;                                                                            // rsp_xbar_demux_011:src0_channel -> rsp_xbar_mux_001:sink11_channel
	wire          rsp_xbar_demux_011_src0_ready;                                                                              // rsp_xbar_mux_001:sink11_ready -> rsp_xbar_demux_011:src0_ready
	wire          rsp_xbar_demux_012_src0_endofpacket;                                                                        // rsp_xbar_demux_012:src0_endofpacket -> rsp_xbar_mux_001:sink12_endofpacket
	wire          rsp_xbar_demux_012_src0_valid;                                                                              // rsp_xbar_demux_012:src0_valid -> rsp_xbar_mux_001:sink12_valid
	wire          rsp_xbar_demux_012_src0_startofpacket;                                                                      // rsp_xbar_demux_012:src0_startofpacket -> rsp_xbar_mux_001:sink12_startofpacket
	wire  [106:0] rsp_xbar_demux_012_src0_data;                                                                               // rsp_xbar_demux_012:src0_data -> rsp_xbar_mux_001:sink12_data
	wire   [15:0] rsp_xbar_demux_012_src0_channel;                                                                            // rsp_xbar_demux_012:src0_channel -> rsp_xbar_mux_001:sink12_channel
	wire          rsp_xbar_demux_012_src0_ready;                                                                              // rsp_xbar_mux_001:sink12_ready -> rsp_xbar_demux_012:src0_ready
	wire          rsp_xbar_demux_014_src0_endofpacket;                                                                        // rsp_xbar_demux_014:src0_endofpacket -> rsp_xbar_mux_001:sink14_endofpacket
	wire          rsp_xbar_demux_014_src0_valid;                                                                              // rsp_xbar_demux_014:src0_valid -> rsp_xbar_mux_001:sink14_valid
	wire          rsp_xbar_demux_014_src0_startofpacket;                                                                      // rsp_xbar_demux_014:src0_startofpacket -> rsp_xbar_mux_001:sink14_startofpacket
	wire  [106:0] rsp_xbar_demux_014_src0_data;                                                                               // rsp_xbar_demux_014:src0_data -> rsp_xbar_mux_001:sink14_data
	wire   [15:0] rsp_xbar_demux_014_src0_channel;                                                                            // rsp_xbar_demux_014:src0_channel -> rsp_xbar_mux_001:sink14_channel
	wire          rsp_xbar_demux_014_src0_ready;                                                                              // rsp_xbar_mux_001:sink14_ready -> rsp_xbar_demux_014:src0_ready
	wire          rsp_xbar_demux_015_src0_endofpacket;                                                                        // rsp_xbar_demux_015:src0_endofpacket -> rsp_xbar_mux_001:sink15_endofpacket
	wire          rsp_xbar_demux_015_src0_valid;                                                                              // rsp_xbar_demux_015:src0_valid -> rsp_xbar_mux_001:sink15_valid
	wire          rsp_xbar_demux_015_src0_startofpacket;                                                                      // rsp_xbar_demux_015:src0_startofpacket -> rsp_xbar_mux_001:sink15_startofpacket
	wire  [106:0] rsp_xbar_demux_015_src0_data;                                                                               // rsp_xbar_demux_015:src0_data -> rsp_xbar_mux_001:sink15_data
	wire   [15:0] rsp_xbar_demux_015_src0_channel;                                                                            // rsp_xbar_demux_015:src0_channel -> rsp_xbar_mux_001:sink15_channel
	wire          rsp_xbar_demux_015_src0_ready;                                                                              // rsp_xbar_mux_001:sink15_ready -> rsp_xbar_demux_015:src0_ready
	wire          addr_router_src_endofpacket;                                                                                // addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          addr_router_src_valid;                                                                                      // addr_router:src_valid -> cmd_xbar_demux:sink_valid
	wire          addr_router_src_startofpacket;                                                                              // addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [106:0] addr_router_src_data;                                                                                       // addr_router:src_data -> cmd_xbar_demux:sink_data
	wire   [15:0] addr_router_src_channel;                                                                                    // addr_router:src_channel -> cmd_xbar_demux:sink_channel
	wire          addr_router_src_ready;                                                                                      // cmd_xbar_demux:sink_ready -> addr_router:src_ready
	wire          rsp_xbar_mux_src_endofpacket;                                                                               // rsp_xbar_mux:src_endofpacket -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_src_valid;                                                                                     // rsp_xbar_mux:src_valid -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_src_startofpacket;                                                                             // rsp_xbar_mux:src_startofpacket -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [106:0] rsp_xbar_mux_src_data;                                                                                      // rsp_xbar_mux:src_data -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [15:0] rsp_xbar_mux_src_channel;                                                                                   // rsp_xbar_mux:src_channel -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_src_ready;                                                                                     // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux:src_ready
	wire          addr_router_001_src_endofpacket;                                                                            // addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire          addr_router_001_src_valid;                                                                                  // addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	wire          addr_router_001_src_startofpacket;                                                                          // addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [106:0] addr_router_001_src_data;                                                                                   // addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	wire   [15:0] addr_router_001_src_channel;                                                                                // addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	wire          addr_router_001_src_ready;                                                                                  // cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	wire          rsp_xbar_mux_001_src_endofpacket;                                                                           // rsp_xbar_mux_001:src_endofpacket -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_001_src_valid;                                                                                 // rsp_xbar_mux_001:src_valid -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_001_src_startofpacket;                                                                         // rsp_xbar_mux_001:src_startofpacket -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [106:0] rsp_xbar_mux_001_src_data;                                                                                  // rsp_xbar_mux_001:src_data -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [15:0] rsp_xbar_mux_001_src_channel;                                                                               // rsp_xbar_mux_001:src_channel -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_001_src_ready;                                                                                 // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_001:src_ready
	wire          addr_router_002_src_endofpacket;                                                                            // addr_router_002:src_endofpacket -> cmd_xbar_demux_002:sink_endofpacket
	wire          addr_router_002_src_valid;                                                                                  // addr_router_002:src_valid -> cmd_xbar_demux_002:sink_valid
	wire          addr_router_002_src_startofpacket;                                                                          // addr_router_002:src_startofpacket -> cmd_xbar_demux_002:sink_startofpacket
	wire   [88:0] addr_router_002_src_data;                                                                                   // addr_router_002:src_data -> cmd_xbar_demux_002:sink_data
	wire   [15:0] addr_router_002_src_channel;                                                                                // addr_router_002:src_channel -> cmd_xbar_demux_002:sink_channel
	wire          addr_router_002_src_ready;                                                                                  // cmd_xbar_demux_002:sink_ready -> addr_router_002:src_ready
	wire          rsp_xbar_demux_010_src1_ready;                                                                              // pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_010:src1_ready
	wire          addr_router_003_src_endofpacket;                                                                            // addr_router_003:src_endofpacket -> cmd_xbar_demux_003:sink_endofpacket
	wire          addr_router_003_src_valid;                                                                                  // addr_router_003:src_valid -> cmd_xbar_demux_003:sink_valid
	wire          addr_router_003_src_startofpacket;                                                                          // addr_router_003:src_startofpacket -> cmd_xbar_demux_003:sink_startofpacket
	wire   [88:0] addr_router_003_src_data;                                                                                   // addr_router_003:src_data -> cmd_xbar_demux_003:sink_data
	wire   [15:0] addr_router_003_src_channel;                                                                                // addr_router_003:src_channel -> cmd_xbar_demux_003:sink_channel
	wire          addr_router_003_src_ready;                                                                                  // cmd_xbar_demux_003:sink_ready -> addr_router_003:src_ready
	wire          rsp_xbar_demux_010_src2_ready;                                                                              // line_drawer_0_avalon_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_010:src2_ready
	wire          cmd_xbar_mux_src_endofpacket;                                                                               // cmd_xbar_mux:src_endofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_src_valid;                                                                                     // cmd_xbar_mux:src_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_src_startofpacket;                                                                             // cmd_xbar_mux:src_startofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_src_data;                                                                                      // cmd_xbar_mux:src_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_mux_src_channel;                                                                                   // cmd_xbar_mux:src_channel -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_src_ready;                                                                                     // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire          id_router_src_endofpacket;                                                                                  // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          id_router_src_valid;                                                                                        // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire          id_router_src_startofpacket;                                                                                // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [106:0] id_router_src_data;                                                                                         // id_router:src_data -> rsp_xbar_demux:sink_data
	wire   [15:0] id_router_src_channel;                                                                                      // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire          id_router_src_ready;                                                                                        // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire          cmd_xbar_mux_001_src_endofpacket;                                                                           // cmd_xbar_mux_001:src_endofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_001_src_valid;                                                                                 // cmd_xbar_mux_001:src_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_001_src_startofpacket;                                                                         // cmd_xbar_mux_001:src_startofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_001_src_data;                                                                                  // cmd_xbar_mux_001:src_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_mux_001_src_channel;                                                                               // cmd_xbar_mux_001:src_channel -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_001_src_ready;                                                                                 // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_001:src_ready
	wire          id_router_001_src_endofpacket;                                                                              // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire          id_router_001_src_valid;                                                                                    // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire          id_router_001_src_startofpacket;                                                                            // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [106:0] id_router_001_src_data;                                                                                     // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire   [15:0] id_router_001_src_channel;                                                                                  // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire          id_router_001_src_ready;                                                                                    // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire          cmd_xbar_mux_002_src_endofpacket;                                                                           // cmd_xbar_mux_002:src_endofpacket -> burst_adapter:sink0_endofpacket
	wire          cmd_xbar_mux_002_src_valid;                                                                                 // cmd_xbar_mux_002:src_valid -> burst_adapter:sink0_valid
	wire          cmd_xbar_mux_002_src_startofpacket;                                                                         // cmd_xbar_mux_002:src_startofpacket -> burst_adapter:sink0_startofpacket
	wire   [88:0] cmd_xbar_mux_002_src_data;                                                                                  // cmd_xbar_mux_002:src_data -> burst_adapter:sink0_data
	wire   [15:0] cmd_xbar_mux_002_src_channel;                                                                               // cmd_xbar_mux_002:src_channel -> burst_adapter:sink0_channel
	wire          cmd_xbar_mux_002_src_ready;                                                                                 // burst_adapter:sink0_ready -> cmd_xbar_mux_002:src_ready
	wire          id_router_002_src_endofpacket;                                                                              // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire          id_router_002_src_valid;                                                                                    // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire          id_router_002_src_startofpacket;                                                                            // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire   [88:0] id_router_002_src_data;                                                                                     // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire   [15:0] id_router_002_src_channel;                                                                                  // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire          id_router_002_src_ready;                                                                                    // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire          cmd_xbar_mux_003_src_endofpacket;                                                                           // cmd_xbar_mux_003:src_endofpacket -> timer_system_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_003_src_valid;                                                                                 // cmd_xbar_mux_003:src_valid -> timer_system_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_003_src_startofpacket;                                                                         // cmd_xbar_mux_003:src_startofpacket -> timer_system_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_003_src_data;                                                                                  // cmd_xbar_mux_003:src_data -> timer_system_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_mux_003_src_channel;                                                                               // cmd_xbar_mux_003:src_channel -> timer_system_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_003_src_ready;                                                                                 // timer_system_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_003:src_ready
	wire          id_router_003_src_endofpacket;                                                                              // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire          id_router_003_src_valid;                                                                                    // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire          id_router_003_src_startofpacket;                                                                            // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [106:0] id_router_003_src_data;                                                                                     // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire   [15:0] id_router_003_src_channel;                                                                                  // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire          id_router_003_src_ready;                                                                                    // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire          cmd_xbar_mux_004_src_endofpacket;                                                                           // cmd_xbar_mux_004:src_endofpacket -> timer_timestamp_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_004_src_valid;                                                                                 // cmd_xbar_mux_004:src_valid -> timer_timestamp_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_004_src_startofpacket;                                                                         // cmd_xbar_mux_004:src_startofpacket -> timer_timestamp_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_004_src_data;                                                                                  // cmd_xbar_mux_004:src_data -> timer_timestamp_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_mux_004_src_channel;                                                                               // cmd_xbar_mux_004:src_channel -> timer_timestamp_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_004_src_ready;                                                                                 // timer_timestamp_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_004:src_ready
	wire          id_router_004_src_endofpacket;                                                                              // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire          id_router_004_src_valid;                                                                                    // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire          id_router_004_src_startofpacket;                                                                            // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [106:0] id_router_004_src_data;                                                                                     // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire   [15:0] id_router_004_src_channel;                                                                                  // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire          id_router_004_src_ready;                                                                                    // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire          cmd_xbar_mux_005_src_endofpacket;                                                                           // cmd_xbar_mux_005:src_endofpacket -> sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_005_src_valid;                                                                                 // cmd_xbar_mux_005:src_valid -> sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_005_src_startofpacket;                                                                         // cmd_xbar_mux_005:src_startofpacket -> sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_005_src_data;                                                                                  // cmd_xbar_mux_005:src_data -> sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_mux_005_src_channel;                                                                               // cmd_xbar_mux_005:src_channel -> sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_005_src_ready;                                                                                 // sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_005:src_ready
	wire          id_router_005_src_endofpacket;                                                                              // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire          id_router_005_src_valid;                                                                                    // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire          id_router_005_src_startofpacket;                                                                            // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [106:0] id_router_005_src_data;                                                                                     // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire   [15:0] id_router_005_src_channel;                                                                                  // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire          id_router_005_src_ready;                                                                                    // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire          cmd_xbar_demux_001_src6_ready;                                                                              // keys_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src6_ready
	wire          id_router_006_src_endofpacket;                                                                              // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire          id_router_006_src_valid;                                                                                    // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire          id_router_006_src_startofpacket;                                                                            // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire  [106:0] id_router_006_src_data;                                                                                     // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire   [15:0] id_router_006_src_channel;                                                                                  // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire          id_router_006_src_ready;                                                                                    // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire          cmd_xbar_demux_001_src7_ready;                                                                              // LEDs_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src7_ready
	wire          id_router_007_src_endofpacket;                                                                              // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire          id_router_007_src_valid;                                                                                    // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire          id_router_007_src_startofpacket;                                                                            // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire  [106:0] id_router_007_src_data;                                                                                     // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire   [15:0] id_router_007_src_channel;                                                                                  // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire          id_router_007_src_ready;                                                                                    // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire          cmd_xbar_demux_001_src8_ready;                                                                              // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src8_ready
	wire          id_router_008_src_endofpacket;                                                                              // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire          id_router_008_src_valid;                                                                                    // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire          id_router_008_src_startofpacket;                                                                            // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire  [106:0] id_router_008_src_data;                                                                                     // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire   [15:0] id_router_008_src_channel;                                                                                  // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire          id_router_008_src_ready;                                                                                    // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire          width_adapter_002_src_ready;                                                                                // burst_adapter_001:sink0_ready -> width_adapter_002:out_ready
	wire          id_router_009_src_endofpacket;                                                                              // id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	wire          id_router_009_src_valid;                                                                                    // id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	wire          id_router_009_src_startofpacket;                                                                            // id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	wire   [79:0] id_router_009_src_data;                                                                                     // id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	wire   [15:0] id_router_009_src_channel;                                                                                  // id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	wire          id_router_009_src_ready;                                                                                    // rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	wire          cmd_xbar_mux_010_src_endofpacket;                                                                           // cmd_xbar_mux_010:src_endofpacket -> burst_adapter_002:sink0_endofpacket
	wire          cmd_xbar_mux_010_src_valid;                                                                                 // cmd_xbar_mux_010:src_valid -> burst_adapter_002:sink0_valid
	wire          cmd_xbar_mux_010_src_startofpacket;                                                                         // cmd_xbar_mux_010:src_startofpacket -> burst_adapter_002:sink0_startofpacket
	wire   [88:0] cmd_xbar_mux_010_src_data;                                                                                  // cmd_xbar_mux_010:src_data -> burst_adapter_002:sink0_data
	wire   [15:0] cmd_xbar_mux_010_src_channel;                                                                               // cmd_xbar_mux_010:src_channel -> burst_adapter_002:sink0_channel
	wire          cmd_xbar_mux_010_src_ready;                                                                                 // burst_adapter_002:sink0_ready -> cmd_xbar_mux_010:src_ready
	wire          id_router_010_src_endofpacket;                                                                              // id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	wire          id_router_010_src_valid;                                                                                    // id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	wire          id_router_010_src_startofpacket;                                                                            // id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	wire   [88:0] id_router_010_src_data;                                                                                     // id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	wire   [15:0] id_router_010_src_channel;                                                                                  // id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	wire          id_router_010_src_ready;                                                                                    // rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	wire          cmd_xbar_demux_001_src11_ready;                                                                             // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src11_ready
	wire          id_router_011_src_endofpacket;                                                                              // id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	wire          id_router_011_src_valid;                                                                                    // id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	wire          id_router_011_src_startofpacket;                                                                            // id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	wire  [106:0] id_router_011_src_data;                                                                                     // id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	wire   [15:0] id_router_011_src_channel;                                                                                  // id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	wire          id_router_011_src_ready;                                                                                    // rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	wire          cmd_xbar_demux_001_src12_ready;                                                                             // line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src12_ready
	wire          id_router_012_src_endofpacket;                                                                              // id_router_012:src_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	wire          id_router_012_src_valid;                                                                                    // id_router_012:src_valid -> rsp_xbar_demux_012:sink_valid
	wire          id_router_012_src_startofpacket;                                                                            // id_router_012:src_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	wire  [106:0] id_router_012_src_data;                                                                                     // id_router_012:src_data -> rsp_xbar_demux_012:sink_data
	wire   [15:0] id_router_012_src_channel;                                                                                  // id_router_012:src_channel -> rsp_xbar_demux_012:sink_channel
	wire          id_router_012_src_ready;                                                                                    // rsp_xbar_demux_012:sink_ready -> id_router_012:src_ready
	wire          width_adapter_004_src_ready;                                                                                // burst_adapter_003:sink0_ready -> width_adapter_004:out_ready
	wire          id_router_013_src_endofpacket;                                                                              // id_router_013:src_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	wire          id_router_013_src_valid;                                                                                    // id_router_013:src_valid -> rsp_xbar_demux_013:sink_valid
	wire          id_router_013_src_startofpacket;                                                                            // id_router_013:src_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	wire   [79:0] id_router_013_src_data;                                                                                     // id_router_013:src_data -> rsp_xbar_demux_013:sink_data
	wire   [15:0] id_router_013_src_channel;                                                                                  // id_router_013:src_channel -> rsp_xbar_demux_013:sink_channel
	wire          id_router_013_src_ready;                                                                                    // rsp_xbar_demux_013:sink_ready -> id_router_013:src_ready
	wire          cmd_xbar_demux_001_src14_ready;                                                                             // pi_request_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src14_ready
	wire          id_router_014_src_endofpacket;                                                                              // id_router_014:src_endofpacket -> rsp_xbar_demux_014:sink_endofpacket
	wire          id_router_014_src_valid;                                                                                    // id_router_014:src_valid -> rsp_xbar_demux_014:sink_valid
	wire          id_router_014_src_startofpacket;                                                                            // id_router_014:src_startofpacket -> rsp_xbar_demux_014:sink_startofpacket
	wire  [106:0] id_router_014_src_data;                                                                                     // id_router_014:src_data -> rsp_xbar_demux_014:sink_data
	wire   [15:0] id_router_014_src_channel;                                                                                  // id_router_014:src_channel -> rsp_xbar_demux_014:sink_channel
	wire          id_router_014_src_ready;                                                                                    // rsp_xbar_demux_014:sink_ready -> id_router_014:src_ready
	wire          cmd_xbar_demux_001_src15_ready;                                                                             // de2_ack_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src15_ready
	wire          id_router_015_src_endofpacket;                                                                              // id_router_015:src_endofpacket -> rsp_xbar_demux_015:sink_endofpacket
	wire          id_router_015_src_valid;                                                                                    // id_router_015:src_valid -> rsp_xbar_demux_015:sink_valid
	wire          id_router_015_src_startofpacket;                                                                            // id_router_015:src_startofpacket -> rsp_xbar_demux_015:sink_startofpacket
	wire  [106:0] id_router_015_src_data;                                                                                     // id_router_015:src_data -> rsp_xbar_demux_015:sink_data
	wire   [15:0] id_router_015_src_channel;                                                                                  // id_router_015:src_channel -> rsp_xbar_demux_015:sink_channel
	wire          id_router_015_src_ready;                                                                                    // rsp_xbar_demux_015:sink_ready -> id_router_015:src_ready
	wire          cmd_xbar_demux_src2_endofpacket;                                                                            // cmd_xbar_demux:src2_endofpacket -> width_adapter:in_endofpacket
	wire          cmd_xbar_demux_src2_valid;                                                                                  // cmd_xbar_demux:src2_valid -> width_adapter:in_valid
	wire          cmd_xbar_demux_src2_startofpacket;                                                                          // cmd_xbar_demux:src2_startofpacket -> width_adapter:in_startofpacket
	wire  [106:0] cmd_xbar_demux_src2_data;                                                                                   // cmd_xbar_demux:src2_data -> width_adapter:in_data
	wire   [15:0] cmd_xbar_demux_src2_channel;                                                                                // cmd_xbar_demux:src2_channel -> width_adapter:in_channel
	wire          cmd_xbar_demux_src2_ready;                                                                                  // width_adapter:in_ready -> cmd_xbar_demux:src2_ready
	wire          width_adapter_src_endofpacket;                                                                              // width_adapter:out_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	wire          width_adapter_src_valid;                                                                                    // width_adapter:out_valid -> cmd_xbar_mux_002:sink0_valid
	wire          width_adapter_src_startofpacket;                                                                            // width_adapter:out_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	wire   [88:0] width_adapter_src_data;                                                                                     // width_adapter:out_data -> cmd_xbar_mux_002:sink0_data
	wire          width_adapter_src_ready;                                                                                    // cmd_xbar_mux_002:sink0_ready -> width_adapter:out_ready
	wire   [15:0] width_adapter_src_channel;                                                                                  // width_adapter:out_channel -> cmd_xbar_mux_002:sink0_channel
	wire          cmd_xbar_demux_001_src2_endofpacket;                                                                        // cmd_xbar_demux_001:src2_endofpacket -> width_adapter_001:in_endofpacket
	wire          cmd_xbar_demux_001_src2_valid;                                                                              // cmd_xbar_demux_001:src2_valid -> width_adapter_001:in_valid
	wire          cmd_xbar_demux_001_src2_startofpacket;                                                                      // cmd_xbar_demux_001:src2_startofpacket -> width_adapter_001:in_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src2_data;                                                                               // cmd_xbar_demux_001:src2_data -> width_adapter_001:in_data
	wire   [15:0] cmd_xbar_demux_001_src2_channel;                                                                            // cmd_xbar_demux_001:src2_channel -> width_adapter_001:in_channel
	wire          cmd_xbar_demux_001_src2_ready;                                                                              // width_adapter_001:in_ready -> cmd_xbar_demux_001:src2_ready
	wire          width_adapter_001_src_endofpacket;                                                                          // width_adapter_001:out_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	wire          width_adapter_001_src_valid;                                                                                // width_adapter_001:out_valid -> cmd_xbar_mux_002:sink1_valid
	wire          width_adapter_001_src_startofpacket;                                                                        // width_adapter_001:out_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	wire   [88:0] width_adapter_001_src_data;                                                                                 // width_adapter_001:out_data -> cmd_xbar_mux_002:sink1_data
	wire          width_adapter_001_src_ready;                                                                                // cmd_xbar_mux_002:sink1_ready -> width_adapter_001:out_ready
	wire   [15:0] width_adapter_001_src_channel;                                                                              // width_adapter_001:out_channel -> cmd_xbar_mux_002:sink1_channel
	wire          cmd_xbar_demux_001_src9_endofpacket;                                                                        // cmd_xbar_demux_001:src9_endofpacket -> width_adapter_002:in_endofpacket
	wire          cmd_xbar_demux_001_src9_valid;                                                                              // cmd_xbar_demux_001:src9_valid -> width_adapter_002:in_valid
	wire          cmd_xbar_demux_001_src9_startofpacket;                                                                      // cmd_xbar_demux_001:src9_startofpacket -> width_adapter_002:in_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src9_data;                                                                               // cmd_xbar_demux_001:src9_data -> width_adapter_002:in_data
	wire   [15:0] cmd_xbar_demux_001_src9_channel;                                                                            // cmd_xbar_demux_001:src9_channel -> width_adapter_002:in_channel
	wire          cmd_xbar_demux_001_src9_ready;                                                                              // width_adapter_002:in_ready -> cmd_xbar_demux_001:src9_ready
	wire          width_adapter_002_src_endofpacket;                                                                          // width_adapter_002:out_endofpacket -> burst_adapter_001:sink0_endofpacket
	wire          width_adapter_002_src_valid;                                                                                // width_adapter_002:out_valid -> burst_adapter_001:sink0_valid
	wire          width_adapter_002_src_startofpacket;                                                                        // width_adapter_002:out_startofpacket -> burst_adapter_001:sink0_startofpacket
	wire   [79:0] width_adapter_002_src_data;                                                                                 // width_adapter_002:out_data -> burst_adapter_001:sink0_data
	wire   [15:0] width_adapter_002_src_channel;                                                                              // width_adapter_002:out_channel -> burst_adapter_001:sink0_channel
	wire          cmd_xbar_demux_001_src10_endofpacket;                                                                       // cmd_xbar_demux_001:src10_endofpacket -> width_adapter_003:in_endofpacket
	wire          cmd_xbar_demux_001_src10_valid;                                                                             // cmd_xbar_demux_001:src10_valid -> width_adapter_003:in_valid
	wire          cmd_xbar_demux_001_src10_startofpacket;                                                                     // cmd_xbar_demux_001:src10_startofpacket -> width_adapter_003:in_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src10_data;                                                                              // cmd_xbar_demux_001:src10_data -> width_adapter_003:in_data
	wire   [15:0] cmd_xbar_demux_001_src10_channel;                                                                           // cmd_xbar_demux_001:src10_channel -> width_adapter_003:in_channel
	wire          cmd_xbar_demux_001_src10_ready;                                                                             // width_adapter_003:in_ready -> cmd_xbar_demux_001:src10_ready
	wire          width_adapter_003_src_endofpacket;                                                                          // width_adapter_003:out_endofpacket -> cmd_xbar_mux_010:sink0_endofpacket
	wire          width_adapter_003_src_valid;                                                                                // width_adapter_003:out_valid -> cmd_xbar_mux_010:sink0_valid
	wire          width_adapter_003_src_startofpacket;                                                                        // width_adapter_003:out_startofpacket -> cmd_xbar_mux_010:sink0_startofpacket
	wire   [88:0] width_adapter_003_src_data;                                                                                 // width_adapter_003:out_data -> cmd_xbar_mux_010:sink0_data
	wire          width_adapter_003_src_ready;                                                                                // cmd_xbar_mux_010:sink0_ready -> width_adapter_003:out_ready
	wire   [15:0] width_adapter_003_src_channel;                                                                              // width_adapter_003:out_channel -> cmd_xbar_mux_010:sink0_channel
	wire          cmd_xbar_demux_001_src13_endofpacket;                                                                       // cmd_xbar_demux_001:src13_endofpacket -> width_adapter_004:in_endofpacket
	wire          cmd_xbar_demux_001_src13_valid;                                                                             // cmd_xbar_demux_001:src13_valid -> width_adapter_004:in_valid
	wire          cmd_xbar_demux_001_src13_startofpacket;                                                                     // cmd_xbar_demux_001:src13_startofpacket -> width_adapter_004:in_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src13_data;                                                                              // cmd_xbar_demux_001:src13_data -> width_adapter_004:in_data
	wire   [15:0] cmd_xbar_demux_001_src13_channel;                                                                           // cmd_xbar_demux_001:src13_channel -> width_adapter_004:in_channel
	wire          cmd_xbar_demux_001_src13_ready;                                                                             // width_adapter_004:in_ready -> cmd_xbar_demux_001:src13_ready
	wire          width_adapter_004_src_endofpacket;                                                                          // width_adapter_004:out_endofpacket -> burst_adapter_003:sink0_endofpacket
	wire          width_adapter_004_src_valid;                                                                                // width_adapter_004:out_valid -> burst_adapter_003:sink0_valid
	wire          width_adapter_004_src_startofpacket;                                                                        // width_adapter_004:out_startofpacket -> burst_adapter_003:sink0_startofpacket
	wire   [79:0] width_adapter_004_src_data;                                                                                 // width_adapter_004:out_data -> burst_adapter_003:sink0_data
	wire   [15:0] width_adapter_004_src_channel;                                                                              // width_adapter_004:out_channel -> burst_adapter_003:sink0_channel
	wire          rsp_xbar_demux_002_src0_endofpacket;                                                                        // rsp_xbar_demux_002:src0_endofpacket -> width_adapter_005:in_endofpacket
	wire          rsp_xbar_demux_002_src0_valid;                                                                              // rsp_xbar_demux_002:src0_valid -> width_adapter_005:in_valid
	wire          rsp_xbar_demux_002_src0_startofpacket;                                                                      // rsp_xbar_demux_002:src0_startofpacket -> width_adapter_005:in_startofpacket
	wire   [88:0] rsp_xbar_demux_002_src0_data;                                                                               // rsp_xbar_demux_002:src0_data -> width_adapter_005:in_data
	wire   [15:0] rsp_xbar_demux_002_src0_channel;                                                                            // rsp_xbar_demux_002:src0_channel -> width_adapter_005:in_channel
	wire          rsp_xbar_demux_002_src0_ready;                                                                              // width_adapter_005:in_ready -> rsp_xbar_demux_002:src0_ready
	wire          width_adapter_005_src_endofpacket;                                                                          // width_adapter_005:out_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire          width_adapter_005_src_valid;                                                                                // width_adapter_005:out_valid -> rsp_xbar_mux:sink2_valid
	wire          width_adapter_005_src_startofpacket;                                                                        // width_adapter_005:out_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [106:0] width_adapter_005_src_data;                                                                                 // width_adapter_005:out_data -> rsp_xbar_mux:sink2_data
	wire          width_adapter_005_src_ready;                                                                                // rsp_xbar_mux:sink2_ready -> width_adapter_005:out_ready
	wire   [15:0] width_adapter_005_src_channel;                                                                              // width_adapter_005:out_channel -> rsp_xbar_mux:sink2_channel
	wire          rsp_xbar_demux_002_src1_endofpacket;                                                                        // rsp_xbar_demux_002:src1_endofpacket -> width_adapter_006:in_endofpacket
	wire          rsp_xbar_demux_002_src1_valid;                                                                              // rsp_xbar_demux_002:src1_valid -> width_adapter_006:in_valid
	wire          rsp_xbar_demux_002_src1_startofpacket;                                                                      // rsp_xbar_demux_002:src1_startofpacket -> width_adapter_006:in_startofpacket
	wire   [88:0] rsp_xbar_demux_002_src1_data;                                                                               // rsp_xbar_demux_002:src1_data -> width_adapter_006:in_data
	wire   [15:0] rsp_xbar_demux_002_src1_channel;                                                                            // rsp_xbar_demux_002:src1_channel -> width_adapter_006:in_channel
	wire          rsp_xbar_demux_002_src1_ready;                                                                              // width_adapter_006:in_ready -> rsp_xbar_demux_002:src1_ready
	wire          width_adapter_006_src_endofpacket;                                                                          // width_adapter_006:out_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire          width_adapter_006_src_valid;                                                                                // width_adapter_006:out_valid -> rsp_xbar_mux_001:sink2_valid
	wire          width_adapter_006_src_startofpacket;                                                                        // width_adapter_006:out_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [106:0] width_adapter_006_src_data;                                                                                 // width_adapter_006:out_data -> rsp_xbar_mux_001:sink2_data
	wire          width_adapter_006_src_ready;                                                                                // rsp_xbar_mux_001:sink2_ready -> width_adapter_006:out_ready
	wire   [15:0] width_adapter_006_src_channel;                                                                              // width_adapter_006:out_channel -> rsp_xbar_mux_001:sink2_channel
	wire          rsp_xbar_demux_009_src0_endofpacket;                                                                        // rsp_xbar_demux_009:src0_endofpacket -> width_adapter_007:in_endofpacket
	wire          rsp_xbar_demux_009_src0_valid;                                                                              // rsp_xbar_demux_009:src0_valid -> width_adapter_007:in_valid
	wire          rsp_xbar_demux_009_src0_startofpacket;                                                                      // rsp_xbar_demux_009:src0_startofpacket -> width_adapter_007:in_startofpacket
	wire   [79:0] rsp_xbar_demux_009_src0_data;                                                                               // rsp_xbar_demux_009:src0_data -> width_adapter_007:in_data
	wire   [15:0] rsp_xbar_demux_009_src0_channel;                                                                            // rsp_xbar_demux_009:src0_channel -> width_adapter_007:in_channel
	wire          rsp_xbar_demux_009_src0_ready;                                                                              // width_adapter_007:in_ready -> rsp_xbar_demux_009:src0_ready
	wire          width_adapter_007_src_endofpacket;                                                                          // width_adapter_007:out_endofpacket -> rsp_xbar_mux_001:sink9_endofpacket
	wire          width_adapter_007_src_valid;                                                                                // width_adapter_007:out_valid -> rsp_xbar_mux_001:sink9_valid
	wire          width_adapter_007_src_startofpacket;                                                                        // width_adapter_007:out_startofpacket -> rsp_xbar_mux_001:sink9_startofpacket
	wire  [106:0] width_adapter_007_src_data;                                                                                 // width_adapter_007:out_data -> rsp_xbar_mux_001:sink9_data
	wire          width_adapter_007_src_ready;                                                                                // rsp_xbar_mux_001:sink9_ready -> width_adapter_007:out_ready
	wire   [15:0] width_adapter_007_src_channel;                                                                              // width_adapter_007:out_channel -> rsp_xbar_mux_001:sink9_channel
	wire          rsp_xbar_demux_010_src0_endofpacket;                                                                        // rsp_xbar_demux_010:src0_endofpacket -> width_adapter_008:in_endofpacket
	wire          rsp_xbar_demux_010_src0_valid;                                                                              // rsp_xbar_demux_010:src0_valid -> width_adapter_008:in_valid
	wire          rsp_xbar_demux_010_src0_startofpacket;                                                                      // rsp_xbar_demux_010:src0_startofpacket -> width_adapter_008:in_startofpacket
	wire   [88:0] rsp_xbar_demux_010_src0_data;                                                                               // rsp_xbar_demux_010:src0_data -> width_adapter_008:in_data
	wire   [15:0] rsp_xbar_demux_010_src0_channel;                                                                            // rsp_xbar_demux_010:src0_channel -> width_adapter_008:in_channel
	wire          rsp_xbar_demux_010_src0_ready;                                                                              // width_adapter_008:in_ready -> rsp_xbar_demux_010:src0_ready
	wire          width_adapter_008_src_endofpacket;                                                                          // width_adapter_008:out_endofpacket -> rsp_xbar_mux_001:sink10_endofpacket
	wire          width_adapter_008_src_valid;                                                                                // width_adapter_008:out_valid -> rsp_xbar_mux_001:sink10_valid
	wire          width_adapter_008_src_startofpacket;                                                                        // width_adapter_008:out_startofpacket -> rsp_xbar_mux_001:sink10_startofpacket
	wire  [106:0] width_adapter_008_src_data;                                                                                 // width_adapter_008:out_data -> rsp_xbar_mux_001:sink10_data
	wire          width_adapter_008_src_ready;                                                                                // rsp_xbar_mux_001:sink10_ready -> width_adapter_008:out_ready
	wire   [15:0] width_adapter_008_src_channel;                                                                              // width_adapter_008:out_channel -> rsp_xbar_mux_001:sink10_channel
	wire          rsp_xbar_demux_013_src0_endofpacket;                                                                        // rsp_xbar_demux_013:src0_endofpacket -> width_adapter_009:in_endofpacket
	wire          rsp_xbar_demux_013_src0_valid;                                                                              // rsp_xbar_demux_013:src0_valid -> width_adapter_009:in_valid
	wire          rsp_xbar_demux_013_src0_startofpacket;                                                                      // rsp_xbar_demux_013:src0_startofpacket -> width_adapter_009:in_startofpacket
	wire   [79:0] rsp_xbar_demux_013_src0_data;                                                                               // rsp_xbar_demux_013:src0_data -> width_adapter_009:in_data
	wire   [15:0] rsp_xbar_demux_013_src0_channel;                                                                            // rsp_xbar_demux_013:src0_channel -> width_adapter_009:in_channel
	wire          rsp_xbar_demux_013_src0_ready;                                                                              // width_adapter_009:in_ready -> rsp_xbar_demux_013:src0_ready
	wire          width_adapter_009_src_endofpacket;                                                                          // width_adapter_009:out_endofpacket -> rsp_xbar_mux_001:sink13_endofpacket
	wire          width_adapter_009_src_valid;                                                                                // width_adapter_009:out_valid -> rsp_xbar_mux_001:sink13_valid
	wire          width_adapter_009_src_startofpacket;                                                                        // width_adapter_009:out_startofpacket -> rsp_xbar_mux_001:sink13_startofpacket
	wire  [106:0] width_adapter_009_src_data;                                                                                 // width_adapter_009:out_data -> rsp_xbar_mux_001:sink13_data
	wire          width_adapter_009_src_ready;                                                                                // rsp_xbar_mux_001:sink13_ready -> width_adapter_009:out_ready
	wire   [15:0] width_adapter_009_src_channel;                                                                              // width_adapter_009:out_channel -> rsp_xbar_mux_001:sink13_channel
	wire          irq_mapper_receiver0_irq;                                                                                   // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire          irq_mapper_receiver1_irq;                                                                                   // timer_system:irq -> irq_mapper:receiver1_irq
	wire          irq_mapper_receiver2_irq;                                                                                   // timer_timestamp:irq -> irq_mapper:receiver2_irq
	wire   [31:0] nios2_qsys_0_d_irq_irq;                                                                                     // irq_mapper:sender_irq -> nios2_qsys_0:d_irq

	nios_system_nios2_qsys_0 nios2_qsys_0 (
		.clk                                   (clocks_sys_clk_clk),                                                        //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                           //                   reset_n.reset_n
		.d_address                             (nios2_qsys_0_data_master_address),                                          //               data_master.address
		.d_byteenable                          (nios2_qsys_0_data_master_byteenable),                                       //                          .byteenable
		.d_read                                (nios2_qsys_0_data_master_read),                                             //                          .read
		.d_readdata                            (nios2_qsys_0_data_master_readdata),                                         //                          .readdata
		.d_waitrequest                         (nios2_qsys_0_data_master_waitrequest),                                      //                          .waitrequest
		.d_write                               (nios2_qsys_0_data_master_write),                                            //                          .write
		.d_writedata                           (nios2_qsys_0_data_master_writedata),                                        //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (nios2_qsys_0_data_master_debugaccess),                                      //                          .debugaccess
		.i_address                             (nios2_qsys_0_instruction_master_address),                                   //        instruction_master.address
		.i_read                                (nios2_qsys_0_instruction_master_read),                                      //                          .read
		.i_readdata                            (nios2_qsys_0_instruction_master_readdata),                                  //                          .readdata
		.i_waitrequest                         (nios2_qsys_0_instruction_master_waitrequest),                               //                          .waitrequest
		.d_irq                                 (nios2_qsys_0_d_irq_irq),                                                    //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_qsys_0_jtag_debug_module_reset_reset),                                //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_read),        //                          .read
		.jtag_debug_module_readdata            (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_write),       //                          .write
		.jtag_debug_module_writedata           (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                                           // custom_instruction_master.readra
	);

	nios_system_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clocks_sys_clk_clk),                                            //   clk1.clk
		.address    (onchip_memory2_0_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.clken      (onchip_memory2_0_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.chipselect (onchip_memory2_0_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.write      (onchip_memory2_0_s1_translator_avalon_anti_slave_0_write),      //       .write
		.readdata   (onchip_memory2_0_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.writedata  (onchip_memory2_0_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (onchip_memory2_0_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                                // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)                             //       .reset_req
	);

	nios_system_keys keys (
		.clk      (clocks_sys_clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address  (keys_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (keys_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (keys_export)                                      // external_connection.export
	);

	nios_system_LEDs leds (
		.clk        (clocks_sys_clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (leds_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~leds_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (leds_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (leds_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (leds_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (leds_export)                                        // external_connection.export
	);

	nios_system_jtag_uart_0 jtag_uart_0 (
		.clk            (clocks_sys_clk_clk),                                                       //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                                          //             reset.reset_n
		.av_chipselect  (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                                  //               irq.irq
	);

	nios_system_sdram sdram (
		.clk            (clocks_sys_clk_clk),                                    //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),                       // reset.reset_n
		.az_addr        (sdram_s1_translator_avalon_anti_slave_0_address),       //    s1.address
		.az_be_n        (~sdram_s1_translator_avalon_anti_slave_0_byteenable),   //      .byteenable_n
		.az_cs          (sdram_s1_translator_avalon_anti_slave_0_chipselect),    //      .chipselect
		.az_data        (sdram_s1_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.az_rd_n        (~sdram_s1_translator_avalon_anti_slave_0_read),         //      .read_n
		.az_wr_n        (~sdram_s1_translator_avalon_anti_slave_0_write),        //      .write_n
		.za_data        (sdram_s1_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.za_valid       (sdram_s1_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.za_waitrequest (sdram_s1_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                                       //  wire.export
		.zs_ba          (sdram_wire_ba),                                         //      .export
		.zs_cas_n       (sdram_wire_cas_n),                                      //      .export
		.zs_cke         (sdram_wire_cke),                                        //      .export
		.zs_cs_n        (sdram_wire_cs_n),                                       //      .export
		.zs_dq          (sdram_wire_dq),                                         //      .export
		.zs_dqm         (sdram_wire_dqm),                                        //      .export
		.zs_ras_n       (sdram_wire_ras_n),                                      //      .export
		.zs_we_n        (sdram_wire_we_n)                                        //      .export
	);

	nios_system_clocks clocks (
		.CLOCK_50    (clk_clk),                            //       clk_in_primary.clk
		.reset       (rst_controller_001_reset_out_reset), // clk_in_primary_reset.reset
		.sys_clk     (clocks_sys_clk_clk),                 //              sys_clk.clk
		.sys_reset_n (),                                   //        sys_clk_reset.reset_n
		.SDRAM_CLK   (sdram_clk_clk),                      //            sdram_clk.clk
		.VGA_CLK     (clocks_vga_clk_clk),                 //              vga_clk.clk
		.CLOCK_27    (clk_27_clk),                         //     clk_in_secondary.clk
		.AUD_CLK     (audio_clk_clk)                       //            audio_clk.clk
	);

	nios_system_character_lcd_0 character_lcd_0 (
		.clk         (clocks_sys_clk_clk),                                                          //        clock_reset.clk
		.reset       (rst_controller_reset_out_reset),                                              //  clock_reset_reset.reset
		.address     (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_address),     //   avalon_lcd_slave.address
		.chipselect  (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_chipselect),  //                   .chipselect
		.read        (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_read),        //                   .read
		.write       (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_write),       //                   .write
		.writedata   (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_writedata),   //                   .writedata
		.readdata    (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_readdata),    //                   .readdata
		.waitrequest (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_waitrequest), //                   .waitrequest
		.LCD_DATA    (lcd_data_DATA),                                                               // external_interface.export
		.LCD_ON      (lcd_data_ON),                                                                 //                   .export
		.LCD_BLON    (lcd_data_BLON),                                                               //                   .export
		.LCD_EN      (lcd_data_EN),                                                                 //                   .export
		.LCD_RS      (lcd_data_RS),                                                                 //                   .export
		.LCD_RW      (lcd_data_RW)                                                                  //                   .export
	);

	nios_system_timer_system timer_system (
		.clk        (clocks_sys_clk_clk),                                        //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                           // reset.reset_n
		.address    (timer_system_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_system_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_system_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_system_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_system_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                                   //   irq.irq
	);

	nios_system_timer_system timer_timestamp (
		.clk        (clocks_sys_clk_clk),                                           //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                              // reset.reset_n
		.address    (timer_timestamp_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_timestamp_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_timestamp_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_timestamp_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_timestamp_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                                      //   irq.irq
	);

	Altera_UP_SD_Card_Avalon_Interface sd_card (
		.i_avalon_chip_select (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_sdcard_slave.chipselect
		.i_avalon_address     (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_address),     //                    .address
		.i_avalon_read        (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_read),        //                    .read
		.i_avalon_write       (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_write),       //                    .write
		.i_avalon_byteenable  (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_byteenable),  //                    .byteenable
		.i_avalon_writedata   (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_writedata),   //                    .writedata
		.o_avalon_readdata    (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_readdata),    //                    .readdata
		.o_avalon_waitrequest (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_waitrequest), //                    .waitrequest
		.i_clock              (clocks_sys_clk_clk),                                                     //          clock_sink.clk
		.i_reset_n            (~rst_controller_reset_out_reset),                                        //    clock_sink_reset.reset_n
		.b_SD_cmd             (sd_card_b_SD_cmd),                                                       //         conduit_end.export
		.b_SD_dat             (sd_card_b_SD_dat),                                                       //                    .export
		.b_SD_dat3            (sd_card_b_SD_dat3),                                                      //                    .export
		.o_SD_clock           (sd_card_o_SD_clock)                                                      //                    .export
	);

	nios_system_pixel_buffer pixel_buffer (
		.clk           (clocks_sys_clk_clk),                                                          //        clock_reset.clk
		.reset         (rst_controller_reset_out_reset),                                              //  clock_reset_reset.reset
		.SRAM_DQ       (sram_pixel_DQ),                                                               // external_interface.export
		.SRAM_ADDR     (sram_pixel_ADDR),                                                             //                   .export
		.SRAM_LB_N     (sram_pixel_LB_N),                                                             //                   .export
		.SRAM_UB_N     (sram_pixel_UB_N),                                                             //                   .export
		.SRAM_CE_N     (sram_pixel_CE_N),                                                             //                   .export
		.SRAM_OE_N     (sram_pixel_OE_N),                                                             //                   .export
		.SRAM_WE_N     (sram_pixel_WE_N),                                                             //                   .export
		.address       (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_address),       //  avalon_sram_slave.address
		.byteenable    (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable),    //                   .byteenable
		.read          (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_read),          //                   .read
		.write         (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_write),         //                   .write
		.writedata     (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_writedata),     //                   .writedata
		.readdata      (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_readdata),      //                   .readdata
		.readdatavalid (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid)  //                   .readdatavalid
	);

	nios_system_pixel_buffer_dma pixel_buffer_dma (
		.clk                  (clocks_sys_clk_clk),                                                              //             clock_reset.clk
		.reset                (rst_controller_reset_out_reset),                                                  //       clock_reset_reset.reset
		.master_readdatavalid (pixel_buffer_dma_avalon_pixel_dma_master_readdatavalid),                          // avalon_pixel_dma_master.readdatavalid
		.master_waitrequest   (pixel_buffer_dma_avalon_pixel_dma_master_waitrequest),                            //                        .waitrequest
		.master_address       (pixel_buffer_dma_avalon_pixel_dma_master_address),                                //                        .address
		.master_arbiterlock   (pixel_buffer_dma_avalon_pixel_dma_master_lock),                                   //                        .lock
		.master_read          (pixel_buffer_dma_avalon_pixel_dma_master_read),                                   //                        .read
		.master_readdata      (pixel_buffer_dma_avalon_pixel_dma_master_readdata),                               //                        .readdata
		.slave_address        (pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_address),    //    avalon_control_slave.address
		.slave_byteenable     (pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_byteenable), //                        .byteenable
		.slave_read           (pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_read),       //                        .read
		.slave_write          (pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_write),      //                        .write
		.slave_writedata      (pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_writedata),  //                        .writedata
		.slave_readdata       (pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_readdata),   //                        .readdata
		.stream_ready         (pixel_buffer_dma_avalon_pixel_source_ready),                                      //     avalon_pixel_source.ready
		.stream_startofpacket (pixel_buffer_dma_avalon_pixel_source_startofpacket),                              //                        .startofpacket
		.stream_endofpacket   (pixel_buffer_dma_avalon_pixel_source_endofpacket),                                //                        .endofpacket
		.stream_valid         (pixel_buffer_dma_avalon_pixel_source_valid),                                      //                        .valid
		.stream_data          (pixel_buffer_dma_avalon_pixel_source_data)                                        //                        .data
	);

	nios_system_rgb_sampler rgb_sampler (
		.clk                      (clocks_sys_clk_clk),                                 //       clock_reset.clk
		.reset                    (rst_controller_reset_out_reset),                     // clock_reset_reset.reset
		.stream_in_startofpacket  (pixel_buffer_dma_avalon_pixel_source_startofpacket), //   avalon_rgb_sink.startofpacket
		.stream_in_endofpacket    (pixel_buffer_dma_avalon_pixel_source_endofpacket),   //                  .endofpacket
		.stream_in_valid          (pixel_buffer_dma_avalon_pixel_source_valid),         //                  .valid
		.stream_in_ready          (pixel_buffer_dma_avalon_pixel_source_ready),         //                  .ready
		.stream_in_data           (pixel_buffer_dma_avalon_pixel_source_data),          //                  .data
		.stream_out_ready         (rgb_sampler_avalon_rgb_source_ready),                // avalon_rgb_source.ready
		.stream_out_startofpacket (rgb_sampler_avalon_rgb_source_startofpacket),        //                  .startofpacket
		.stream_out_endofpacket   (rgb_sampler_avalon_rgb_source_endofpacket),          //                  .endofpacket
		.stream_out_valid         (rgb_sampler_avalon_rgb_source_valid),                //                  .valid
		.stream_out_data          (rgb_sampler_avalon_rgb_source_data)                  //                  .data
	);

	nios_system_scaler scaler (
		.clk                      (clocks_sys_clk_clk),                          //          clock_reset.clk
		.reset                    (rst_controller_reset_out_reset),              //    clock_reset_reset.reset
		.stream_in_startofpacket  (rgb_sampler_avalon_rgb_source_startofpacket), //   avalon_scaler_sink.startofpacket
		.stream_in_endofpacket    (rgb_sampler_avalon_rgb_source_endofpacket),   //                     .endofpacket
		.stream_in_valid          (rgb_sampler_avalon_rgb_source_valid),         //                     .valid
		.stream_in_ready          (rgb_sampler_avalon_rgb_source_ready),         //                     .ready
		.stream_in_data           (rgb_sampler_avalon_rgb_source_data),          //                     .data
		.stream_out_ready         (scaler_avalon_scaler_source_ready),           // avalon_scaler_source.ready
		.stream_out_startofpacket (scaler_avalon_scaler_source_startofpacket),   //                     .startofpacket
		.stream_out_endofpacket   (scaler_avalon_scaler_source_endofpacket),     //                     .endofpacket
		.stream_out_valid         (scaler_avalon_scaler_source_valid),           //                     .valid
		.stream_out_data          (scaler_avalon_scaler_source_data)             //                     .data
	);

	nios_system_video_fifo video_fifo (
		.clk_stream_in            (clocks_sys_clk_clk),                               //         clock_stream_in.clk
		.reset_stream_in          (rst_controller_reset_out_reset),                   //   clock_stream_in_reset.reset
		.clk_stream_out           (clocks_vga_clk_clk),                               //        clock_stream_out.clk
		.reset_stream_out         (rst_controller_002_reset_out_reset),               //  clock_stream_out_reset.reset
		.stream_in_ready          (scaler_avalon_scaler_source_ready),                //   avalon_dc_buffer_sink.ready
		.stream_in_startofpacket  (scaler_avalon_scaler_source_startofpacket),        //                        .startofpacket
		.stream_in_endofpacket    (scaler_avalon_scaler_source_endofpacket),          //                        .endofpacket
		.stream_in_valid          (scaler_avalon_scaler_source_valid),                //                        .valid
		.stream_in_data           (scaler_avalon_scaler_source_data),                 //                        .data
		.stream_out_ready         (video_fifo_avalon_dc_buffer_source_ready),         // avalon_dc_buffer_source.ready
		.stream_out_startofpacket (video_fifo_avalon_dc_buffer_source_startofpacket), //                        .startofpacket
		.stream_out_endofpacket   (video_fifo_avalon_dc_buffer_source_endofpacket),   //                        .endofpacket
		.stream_out_valid         (video_fifo_avalon_dc_buffer_source_valid),         //                        .valid
		.stream_out_data          (video_fifo_avalon_dc_buffer_source_data)           //                        .data
	);

	nios_system_vga_controller vga_controller (
		.clk           (clocks_vga_clk_clk),                               //        clock_reset.clk
		.reset         (rst_controller_002_reset_out_reset),               //  clock_reset_reset.reset
		.data          (video_fifo_avalon_dc_buffer_source_data),          //    avalon_vga_sink.data
		.startofpacket (video_fifo_avalon_dc_buffer_source_startofpacket), //                   .startofpacket
		.endofpacket   (video_fifo_avalon_dc_buffer_source_endofpacket),   //                   .endofpacket
		.valid         (video_fifo_avalon_dc_buffer_source_valid),         //                   .valid
		.ready         (video_fifo_avalon_dc_buffer_source_ready),         //                   .ready
		.VGA_CLK       (vga_controller_CLK),                               // external_interface.export
		.VGA_HS        (vga_controller_HS),                                //                   .export
		.VGA_VS        (vga_controller_VS),                                //                   .export
		.VGA_BLANK     (vga_controller_BLANK),                             //                   .export
		.VGA_SYNC      (vga_controller_SYNC),                              //                   .export
		.VGA_R         (vga_controller_R),                                 //                   .export
		.VGA_G         (vga_controller_G),                                 //                   .export
		.VGA_B         (vga_controller_B)                                  //                   .export
	);

	line_drawer line_drawer_0 (
		.clk                (clocks_sys_clk_clk),                                                    //          clock.clk
		.reset_n            (~rst_controller_reset_out_reset),                                       //          reset.reset_n
		.slave_addr         (line_drawer_0_avalon_slave_0_translator_avalon_anti_slave_0_address),   // avalon_slave_0.address
		.slave_rd_en        (line_drawer_0_avalon_slave_0_translator_avalon_anti_slave_0_read),      //               .read
		.slave_wr_en        (line_drawer_0_avalon_slave_0_translator_avalon_anti_slave_0_write),     //               .write
		.slave_readdata     (line_drawer_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),  //               .readdata
		.slave_writedata    (line_drawer_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata), //               .writedata
		.master_rd_en       (line_drawer_0_avalon_master_read),                                      //  avalon_master.read
		.master_wr_en       (line_drawer_0_avalon_master_write),                                     //               .write
		.master_be          (line_drawer_0_avalon_master_byteenable),                                //               .byteenable
		.master_readdata    (line_drawer_0_avalon_master_readdata),                                  //               .readdata
		.master_writedata   (line_drawer_0_avalon_master_writedata),                                 //               .writedata
		.master_waitrequest (line_drawer_0_avalon_master_waitrequest),                               //               .waitrequest
		.master_addr        (line_drawer_0_avalon_master_address)                                    //               .address
	);

	nios_system_dual_port_ram dual_port_ram (
		.clk         (clocks_sys_clk_clk),                                         //   clk1.clk
		.address     (dual_port_ram_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.clken       (dual_port_ram_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.chipselect  (dual_port_ram_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.write       (dual_port_ram_s1_translator_avalon_anti_slave_0_write),      //       .write
		.readdata    (dual_port_ram_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.writedata   (dual_port_ram_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.reset       (rst_controller_reset_out_reset),                             // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),                         //       .reset_req
		.address2    (dual_port_ram_s2_address),                                   //     s2.address
		.chipselect2 (dual_port_ram_s2_chipselect),                                //       .chipselect
		.clken2      (dual_port_ram_s2_clken),                                     //       .clken
		.write2      (dual_port_ram_s2_write),                                     //       .write
		.readdata2   (dual_port_ram_s2_readdata),                                  //       .readdata
		.writedata2  (dual_port_ram_s2_writedata),                                 //       .writedata
		.clk2        (clk_pi_clk),                                                 //   clk2.clk
		.reset2      (rst_controller_003_reset_out_reset),                         // reset2.reset
		.reset_req2  (rst_controller_003_reset_out_reset_req)                      //       .reset_req
	);

	nios_system_de2_ack de2_ack (
		.clk        (clocks_sys_clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                      //               reset.reset_n
		.address    (de2_ack_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~de2_ack_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (de2_ack_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (de2_ack_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (de2_ack_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (de2_ack_export)                                        // external_connection.export
	);

	nios_system_pi_request pi_request (
		.clk      (clocks_sys_clk_clk),                                    //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //               reset.reset_n
		.address  (pi_request_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (pi_request_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (pi_request_export)                                      // external_connection.export
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (25),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios2_qsys_0_instruction_master_translator (
		.clk                      (clocks_sys_clk_clk),                                                                 //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                     //                     reset.reset
		.uav_address              (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (nios2_qsys_0_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (nios2_qsys_0_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read                  (nios2_qsys_0_instruction_master_read),                                               //                          .read
		.av_readdata              (nios2_qsys_0_instruction_master_readdata),                                           //                          .readdata
		.av_burstcount            (1'b1),                                                                               //               (terminated)
		.av_byteenable            (4'b1111),                                                                            //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                               //               (terminated)
		.av_begintransfer         (1'b0),                                                                               //               (terminated)
		.av_chipselect            (1'b0),                                                                               //               (terminated)
		.av_readdatavalid         (),                                                                                   //               (terminated)
		.av_write                 (1'b0),                                                                               //               (terminated)
		.av_writedata             (32'b00000000000000000000000000000000),                                               //               (terminated)
		.av_lock                  (1'b0),                                                                               //               (terminated)
		.av_debugaccess           (1'b0),                                                                               //               (terminated)
		.uav_clken                (),                                                                                   //               (terminated)
		.av_clken                 (1'b1),                                                                               //               (terminated)
		.uav_response             (2'b00),                                                                              //               (terminated)
		.av_response              (),                                                                                   //               (terminated)
		.uav_writeresponserequest (),                                                                                   //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                               //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                               //               (terminated)
		.av_writeresponsevalid    ()                                                                                    //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (25),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (1)
	) nios2_qsys_0_data_master_translator (
		.clk                      (clocks_sys_clk_clk),                                                          //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                              //                     reset.reset
		.uav_address              (nios2_qsys_0_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (nios2_qsys_0_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (nios2_qsys_0_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (nios2_qsys_0_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (nios2_qsys_0_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (nios2_qsys_0_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (nios2_qsys_0_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (nios2_qsys_0_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (nios2_qsys_0_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (nios2_qsys_0_data_master_byteenable),                                         //                          .byteenable
		.av_read                  (nios2_qsys_0_data_master_read),                                               //                          .read
		.av_readdata              (nios2_qsys_0_data_master_readdata),                                           //                          .readdata
		.av_write                 (nios2_qsys_0_data_master_write),                                              //                          .write
		.av_writedata             (nios2_qsys_0_data_master_writedata),                                          //                          .writedata
		.av_debugaccess           (nios2_qsys_0_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount            (1'b1),                                                                        //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                        //               (terminated)
		.av_begintransfer         (1'b0),                                                                        //               (terminated)
		.av_chipselect            (1'b0),                                                                        //               (terminated)
		.av_readdatavalid         (),                                                                            //               (terminated)
		.av_lock                  (1'b0),                                                                        //               (terminated)
		.uav_clken                (),                                                                            //               (terminated)
		.av_clken                 (1'b1),                                                                        //               (terminated)
		.uav_response             (2'b00),                                                                       //               (terminated)
		.av_response              (),                                                                            //               (terminated)
		.uav_writeresponserequest (),                                                                            //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                        //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                        //               (terminated)
		.av_writeresponsevalid    ()                                                                             //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (16),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (2),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (2),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (2),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) pixel_buffer_dma_avalon_pixel_dma_master_translator (
		.clk                      (clocks_sys_clk_clk),                                                                          //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                              //                     reset.reset
		.uav_address              (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (pixel_buffer_dma_avalon_pixel_dma_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (pixel_buffer_dma_avalon_pixel_dma_master_waitrequest),                                        //                          .waitrequest
		.av_read                  (pixel_buffer_dma_avalon_pixel_dma_master_read),                                               //                          .read
		.av_readdata              (pixel_buffer_dma_avalon_pixel_dma_master_readdata),                                           //                          .readdata
		.av_readdatavalid         (pixel_buffer_dma_avalon_pixel_dma_master_readdatavalid),                                      //                          .readdatavalid
		.av_lock                  (pixel_buffer_dma_avalon_pixel_dma_master_lock),                                               //                          .lock
		.av_burstcount            (1'b1),                                                                                        //               (terminated)
		.av_byteenable            (2'b11),                                                                                       //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                                        //               (terminated)
		.av_begintransfer         (1'b0),                                                                                        //               (terminated)
		.av_chipselect            (1'b0),                                                                                        //               (terminated)
		.av_write                 (1'b0),                                                                                        //               (terminated)
		.av_writedata             (16'b0000000000000000),                                                                        //               (terminated)
		.av_debugaccess           (1'b0),                                                                                        //               (terminated)
		.uav_clken                (),                                                                                            //               (terminated)
		.av_clken                 (1'b1),                                                                                        //               (terminated)
		.uav_response             (2'b00),                                                                                       //               (terminated)
		.av_response              (),                                                                                            //               (terminated)
		.uav_writeresponserequest (),                                                                                            //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                                        //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                                        //               (terminated)
		.av_writeresponsevalid    ()                                                                                             //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (16),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (2),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (2),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (2),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) line_drawer_0_avalon_master_translator (
		.clk                      (clocks_sys_clk_clk),                                                             //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                 //                     reset.reset
		.uav_address              (line_drawer_0_avalon_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (line_drawer_0_avalon_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (line_drawer_0_avalon_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (line_drawer_0_avalon_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (line_drawer_0_avalon_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (line_drawer_0_avalon_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (line_drawer_0_avalon_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (line_drawer_0_avalon_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (line_drawer_0_avalon_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (line_drawer_0_avalon_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (line_drawer_0_avalon_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (line_drawer_0_avalon_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (line_drawer_0_avalon_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (line_drawer_0_avalon_master_byteenable),                                         //                          .byteenable
		.av_read                  (line_drawer_0_avalon_master_read),                                               //                          .read
		.av_readdata              (line_drawer_0_avalon_master_readdata),                                           //                          .readdata
		.av_write                 (line_drawer_0_avalon_master_write),                                              //                          .write
		.av_writedata             (line_drawer_0_avalon_master_writedata),                                          //                          .writedata
		.av_burstcount            (1'b1),                                                                           //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                           //               (terminated)
		.av_begintransfer         (1'b0),                                                                           //               (terminated)
		.av_chipselect            (1'b0),                                                                           //               (terminated)
		.av_readdatavalid         (),                                                                               //               (terminated)
		.av_lock                  (1'b0),                                                                           //               (terminated)
		.av_debugaccess           (1'b0),                                                                           //               (terminated)
		.uav_clken                (),                                                                               //               (terminated)
		.av_clken                 (1'b1),                                                                           //               (terminated)
		.uav_response             (2'b00),                                                                          //               (terminated)
		.av_response              (),                                                                               //               (terminated)
		.uav_writeresponserequest (),                                                                               //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                           //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                           //               (terminated)
		.av_writeresponsevalid    ()                                                                                //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) nios2_qsys_0_jtag_debug_module_translator (
		.clk                      (clocks_sys_clk_clk),                                                                        //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                            //                    reset.reset
		.uav_address              (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess           (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer         (),                                                                                          //              (terminated)
		.av_beginbursttransfer    (),                                                                                          //              (terminated)
		.av_burstcount            (),                                                                                          //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                      //              (terminated)
		.av_writebyteenable       (),                                                                                          //              (terminated)
		.av_lock                  (),                                                                                          //              (terminated)
		.av_chipselect            (),                                                                                          //              (terminated)
		.av_clken                 (),                                                                                          //              (terminated)
		.uav_clken                (1'b0),                                                                                      //              (terminated)
		.av_outputenable          (),                                                                                          //              (terminated)
		.uav_response             (),                                                                                          //              (terminated)
		.av_response              (2'b00),                                                                                     //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                      //              (terminated)
		.uav_writeresponsevalid   (),                                                                                          //              (terminated)
		.av_writeresponserequest  (),                                                                                          //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (10),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) onchip_memory2_0_s1_translator (
		.clk                      (clocks_sys_clk_clk),                                                             //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                 //                    reset.reset
		.uav_address              (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (onchip_memory2_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (onchip_memory2_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (onchip_memory2_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (onchip_memory2_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (onchip_memory2_0_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (onchip_memory2_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken                 (onchip_memory2_0_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read                  (),                                                                               //              (terminated)
		.av_begintransfer         (),                                                                               //              (terminated)
		.av_beginbursttransfer    (),                                                                               //              (terminated)
		.av_burstcount            (),                                                                               //              (terminated)
		.av_readdatavalid         (1'b0),                                                                           //              (terminated)
		.av_waitrequest           (1'b0),                                                                           //              (terminated)
		.av_writebyteenable       (),                                                                               //              (terminated)
		.av_lock                  (),                                                                               //              (terminated)
		.uav_clken                (1'b0),                                                                           //              (terminated)
		.av_debugaccess           (),                                                                               //              (terminated)
		.av_outputenable          (),                                                                               //              (terminated)
		.uav_response             (),                                                                               //              (terminated)
		.av_response              (2'b00),                                                                          //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                           //              (terminated)
		.uav_writeresponsevalid   (),                                                                               //              (terminated)
		.av_writeresponserequest  (),                                                                               //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                            //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (22),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sdram_s1_translator (
		.clk                      (clocks_sys_clk_clk),                                                  //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                      //                    reset.reset
		.uav_address              (sdram_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sdram_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sdram_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (sdram_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (sdram_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (sdram_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (sdram_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (sdram_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (sdram_s1_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest           (sdram_s1_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (sdram_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                    //              (terminated)
		.av_burstcount            (),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                    //              (terminated)
		.av_lock                  (),                                                                    //              (terminated)
		.av_clken                 (),                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                //              (terminated)
		.av_debugaccess           (),                                                                    //              (terminated)
		.av_outputenable          (),                                                                    //              (terminated)
		.uav_response             (),                                                                    //              (terminated)
		.av_response              (2'b00),                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_system_s1_translator (
		.clk                      (clocks_sys_clk_clk),                                                         //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                             //                    reset.reset
		.uav_address              (timer_system_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (timer_system_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (timer_system_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (timer_system_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (timer_system_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (timer_system_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (timer_system_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (timer_system_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (timer_system_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (timer_system_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (timer_system_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (timer_system_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (timer_system_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (timer_system_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (timer_system_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (timer_system_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                           //              (terminated)
		.av_begintransfer         (),                                                                           //              (terminated)
		.av_beginbursttransfer    (),                                                                           //              (terminated)
		.av_burstcount            (),                                                                           //              (terminated)
		.av_byteenable            (),                                                                           //              (terminated)
		.av_readdatavalid         (1'b0),                                                                       //              (terminated)
		.av_waitrequest           (1'b0),                                                                       //              (terminated)
		.av_writebyteenable       (),                                                                           //              (terminated)
		.av_lock                  (),                                                                           //              (terminated)
		.av_clken                 (),                                                                           //              (terminated)
		.uav_clken                (1'b0),                                                                       //              (terminated)
		.av_debugaccess           (),                                                                           //              (terminated)
		.av_outputenable          (),                                                                           //              (terminated)
		.uav_response             (),                                                                           //              (terminated)
		.av_response              (2'b00),                                                                      //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                       //              (terminated)
		.uav_writeresponsevalid   (),                                                                           //              (terminated)
		.av_writeresponserequest  (),                                                                           //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_timestamp_s1_translator (
		.clk                      (clocks_sys_clk_clk),                                                            //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                //                    reset.reset
		.uav_address              (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (timer_timestamp_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (timer_timestamp_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (timer_timestamp_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (timer_timestamp_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (timer_timestamp_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                              //              (terminated)
		.av_begintransfer         (),                                                                              //              (terminated)
		.av_beginbursttransfer    (),                                                                              //              (terminated)
		.av_burstcount            (),                                                                              //              (terminated)
		.av_byteenable            (),                                                                              //              (terminated)
		.av_readdatavalid         (1'b0),                                                                          //              (terminated)
		.av_waitrequest           (1'b0),                                                                          //              (terminated)
		.av_writebyteenable       (),                                                                              //              (terminated)
		.av_lock                  (),                                                                              //              (terminated)
		.av_clken                 (),                                                                              //              (terminated)
		.uav_clken                (1'b0),                                                                          //              (terminated)
		.av_debugaccess           (),                                                                              //              (terminated)
		.av_outputenable          (),                                                                              //              (terminated)
		.uav_response             (),                                                                              //              (terminated)
		.av_response              (2'b00),                                                                         //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                          //              (terminated)
		.uav_writeresponsevalid   (),                                                                              //              (terminated)
		.av_writeresponserequest  (),                                                                              //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                           //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (8),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sd_card_avalon_sdcard_slave_translator (
		.clk                      (clocks_sys_clk_clk),                                                                     //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                         //                    reset.reset
		.uav_address              (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                                       //              (terminated)
		.av_burstcount            (),                                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                                       //              (terminated)
		.av_lock                  (),                                                                                       //              (terminated)
		.av_clken                 (),                                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                                   //              (terminated)
		.av_debugaccess           (),                                                                                       //              (terminated)
		.av_outputenable          (),                                                                                       //              (terminated)
		.uav_response             (),                                                                                       //              (terminated)
		.av_response              (2'b00),                                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) keys_s1_translator (
		.clk                      (clocks_sys_clk_clk),                                                 //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address              (keys_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (keys_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (keys_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (keys_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (keys_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (keys_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (keys_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (keys_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (keys_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (keys_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (keys_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (keys_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (keys_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                   //              (terminated)
		.av_read                  (),                                                                   //              (terminated)
		.av_writedata             (),                                                                   //              (terminated)
		.av_begintransfer         (),                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                   //              (terminated)
		.av_burstcount            (),                                                                   //              (terminated)
		.av_byteenable            (),                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                               //              (terminated)
		.av_writebyteenable       (),                                                                   //              (terminated)
		.av_lock                  (),                                                                   //              (terminated)
		.av_chipselect            (),                                                                   //              (terminated)
		.av_clken                 (),                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                               //              (terminated)
		.av_debugaccess           (),                                                                   //              (terminated)
		.av_outputenable          (),                                                                   //              (terminated)
		.uav_response             (),                                                                   //              (terminated)
		.av_response              (2'b00),                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) leds_s1_translator (
		.clk                      (clocks_sys_clk_clk),                                                 //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address              (leds_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (leds_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (leds_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (leds_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (leds_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (leds_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (leds_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (leds_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (leds_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (leds_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (leds_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (leds_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (leds_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (leds_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (leds_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (leds_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                   //              (terminated)
		.av_begintransfer         (),                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                   //              (terminated)
		.av_burstcount            (),                                                                   //              (terminated)
		.av_byteenable            (),                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                               //              (terminated)
		.av_writebyteenable       (),                                                                   //              (terminated)
		.av_lock                  (),                                                                   //              (terminated)
		.av_clken                 (),                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                               //              (terminated)
		.av_debugaccess           (),                                                                   //              (terminated)
		.av_outputenable          (),                                                                   //              (terminated)
		.uav_response             (),                                                                   //              (terminated)
		.av_response              (2'b00),                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_0_avalon_jtag_slave_translator (
		.clk                      (clocks_sys_clk_clk),                                                                       //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                           //                    reset.reset
		.uav_address              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                                         //              (terminated)
		.av_burstcount            (),                                                                                         //              (terminated)
		.av_byteenable            (),                                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                                         //              (terminated)
		.av_lock                  (),                                                                                         //              (terminated)
		.av_clken                 (),                                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                                     //              (terminated)
		.av_debugaccess           (),                                                                                         //              (terminated)
		.av_outputenable          (),                                                                                         //              (terminated)
		.uav_response             (),                                                                                         //              (terminated)
		.av_response              (2'b00),                                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) character_lcd_0_avalon_lcd_slave_translator (
		.clk                      (clocks_sys_clk_clk),                                                                          //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                              //                    reset.reset
		.uav_address              (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                            //              (terminated)
		.av_beginbursttransfer    (),                                                                                            //              (terminated)
		.av_burstcount            (),                                                                                            //              (terminated)
		.av_byteenable            (),                                                                                            //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                        //              (terminated)
		.av_writebyteenable       (),                                                                                            //              (terminated)
		.av_lock                  (),                                                                                            //              (terminated)
		.av_clken                 (),                                                                                            //              (terminated)
		.uav_clken                (1'b0),                                                                                        //              (terminated)
		.av_debugaccess           (),                                                                                            //              (terminated)
		.av_outputenable          (),                                                                                            //              (terminated)
		.uav_response             (),                                                                                            //              (terminated)
		.av_response              (2'b00),                                                                                       //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                        //              (terminated)
		.uav_writeresponsevalid   (),                                                                                            //              (terminated)
		.av_writeresponserequest  (),                                                                                            //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (18),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pixel_buffer_avalon_sram_slave_translator (
		.clk                      (clocks_sys_clk_clk),                                                                        //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                            //                    reset.reset
		.uav_address              (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_begintransfer         (),                                                                                          //              (terminated)
		.av_beginbursttransfer    (),                                                                                          //              (terminated)
		.av_burstcount            (),                                                                                          //              (terminated)
		.av_waitrequest           (1'b0),                                                                                      //              (terminated)
		.av_writebyteenable       (),                                                                                          //              (terminated)
		.av_lock                  (),                                                                                          //              (terminated)
		.av_chipselect            (),                                                                                          //              (terminated)
		.av_clken                 (),                                                                                          //              (terminated)
		.uav_clken                (1'b0),                                                                                      //              (terminated)
		.av_debugaccess           (),                                                                                          //              (terminated)
		.av_outputenable          (),                                                                                          //              (terminated)
		.uav_response             (),                                                                                          //              (terminated)
		.av_response              (2'b00),                                                                                     //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                      //              (terminated)
		.uav_writeresponsevalid   (),                                                                                          //              (terminated)
		.av_writeresponserequest  (),                                                                                          //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pixel_buffer_dma_avalon_control_slave_translator (
		.clk                      (clocks_sys_clk_clk),                                                                               //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                                   //                    reset.reset
		.uav_address              (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_begintransfer         (),                                                                                                 //              (terminated)
		.av_beginbursttransfer    (),                                                                                                 //              (terminated)
		.av_burstcount            (),                                                                                                 //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                             //              (terminated)
		.av_waitrequest           (1'b0),                                                                                             //              (terminated)
		.av_writebyteenable       (),                                                                                                 //              (terminated)
		.av_lock                  (),                                                                                                 //              (terminated)
		.av_chipselect            (),                                                                                                 //              (terminated)
		.av_clken                 (),                                                                                                 //              (terminated)
		.uav_clken                (1'b0),                                                                                             //              (terminated)
		.av_debugaccess           (),                                                                                                 //              (terminated)
		.av_outputenable          (),                                                                                                 //              (terminated)
		.uav_response             (),                                                                                                 //              (terminated)
		.av_response              (2'b00),                                                                                            //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                             //              (terminated)
		.uav_writeresponsevalid   (),                                                                                                 //              (terminated)
		.av_writeresponserequest  (),                                                                                                 //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) line_drawer_0_avalon_slave_0_translator (
		.clk                      (clocks_sys_clk_clk),                                                                      //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                          //                    reset.reset
		.uav_address              (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (line_drawer_0_avalon_slave_0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (line_drawer_0_avalon_slave_0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (line_drawer_0_avalon_slave_0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (line_drawer_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (line_drawer_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer         (),                                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                                        //              (terminated)
		.av_burstcount            (),                                                                                        //              (terminated)
		.av_byteenable            (),                                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                                        //              (terminated)
		.av_lock                  (),                                                                                        //              (terminated)
		.av_chipselect            (),                                                                                        //              (terminated)
		.av_clken                 (),                                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                                    //              (terminated)
		.av_debugaccess           (),                                                                                        //              (terminated)
		.av_outputenable          (),                                                                                        //              (terminated)
		.uav_response             (),                                                                                        //              (terminated)
		.av_response              (2'b00),                                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (12),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) dual_port_ram_s1_translator (
		.clk                      (clocks_sys_clk_clk),                                                          //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                              //                    reset.reset
		.uav_address              (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (dual_port_ram_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (dual_port_ram_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (dual_port_ram_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (dual_port_ram_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (dual_port_ram_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken                 (dual_port_ram_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read                  (),                                                                            //              (terminated)
		.av_begintransfer         (),                                                                            //              (terminated)
		.av_beginbursttransfer    (),                                                                            //              (terminated)
		.av_burstcount            (),                                                                            //              (terminated)
		.av_byteenable            (),                                                                            //              (terminated)
		.av_readdatavalid         (1'b0),                                                                        //              (terminated)
		.av_waitrequest           (1'b0),                                                                        //              (terminated)
		.av_writebyteenable       (),                                                                            //              (terminated)
		.av_lock                  (),                                                                            //              (terminated)
		.uav_clken                (1'b0),                                                                        //              (terminated)
		.av_debugaccess           (),                                                                            //              (terminated)
		.av_outputenable          (),                                                                            //              (terminated)
		.uav_response             (),                                                                            //              (terminated)
		.av_response              (2'b00),                                                                       //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                        //              (terminated)
		.uav_writeresponsevalid   (),                                                                            //              (terminated)
		.av_writeresponserequest  (),                                                                            //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pi_request_s1_translator (
		.clk                      (clocks_sys_clk_clk),                                                       //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                           //                    reset.reset
		.uav_address              (pi_request_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (pi_request_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (pi_request_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (pi_request_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (pi_request_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (pi_request_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (pi_request_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (pi_request_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (pi_request_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (pi_request_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (pi_request_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (pi_request_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (pi_request_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                         //              (terminated)
		.av_read                  (),                                                                         //              (terminated)
		.av_writedata             (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_chipselect            (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) de2_ack_s1_translator (
		.clk                      (clocks_sys_clk_clk),                                                    //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address              (de2_ack_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (de2_ack_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (de2_ack_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (de2_ack_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (de2_ack_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (de2_ack_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (de2_ack_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (de2_ack_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (de2_ack_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (de2_ack_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (de2_ack_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (de2_ack_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (de2_ack_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (de2_ack_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (de2_ack_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (de2_ack_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                      //              (terminated)
		.av_begintransfer         (),                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                      //              (terminated)
		.av_burstcount            (),                                                                      //              (terminated)
		.av_byteenable            (),                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                      //              (terminated)
		.av_lock                  (),                                                                      //              (terminated)
		.av_clken                 (),                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                  //              (terminated)
		.av_debugaccess           (),                                                                      //              (terminated)
		.av_outputenable          (),                                                                      //              (terminated)
		.uav_response             (),                                                                      //              (terminated)
		.av_response              (2'b00),                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                   //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_BEGIN_BURST           (87),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_THREAD_ID_H           (97),
		.PKT_THREAD_ID_L           (97),
		.PKT_CACHE_H               (104),
		.PKT_CACHE_L               (101),
		.PKT_DATA_SIDEBAND_H       (86),
		.PKT_DATA_SIDEBAND_L       (86),
		.PKT_QOS_H                 (88),
		.PKT_QOS_L                 (88),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (16),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (2),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                          //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.av_address              (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_mux_src_valid),                                                                      //        rp.valid
		.rp_data                 (rsp_xbar_mux_src_data),                                                                       //          .data
		.rp_channel              (rsp_xbar_mux_src_channel),                                                                    //          .channel
		.rp_startofpacket        (rsp_xbar_mux_src_startofpacket),                                                              //          .startofpacket
		.rp_endofpacket          (rsp_xbar_mux_src_endofpacket),                                                                //          .endofpacket
		.rp_ready                (rsp_xbar_mux_src_ready),                                                                      //          .ready
		.av_response             (),                                                                                            // (terminated)
		.av_writeresponserequest (1'b0),                                                                                        // (terminated)
		.av_writeresponsevalid   ()                                                                                             // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_BEGIN_BURST           (87),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_THREAD_ID_H           (97),
		.PKT_THREAD_ID_L           (97),
		.PKT_CACHE_H               (104),
		.PKT_CACHE_L               (101),
		.PKT_DATA_SIDEBAND_H       (86),
		.PKT_DATA_SIDEBAND_L       (86),
		.PKT_QOS_H                 (88),
		.PKT_QOS_L                 (88),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (16),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                   //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.av_address              (nios2_qsys_0_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (nios2_qsys_0_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (nios2_qsys_0_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (nios2_qsys_0_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (nios2_qsys_0_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (nios2_qsys_0_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (nios2_qsys_0_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_mux_001_src_valid),                                                           //        rp.valid
		.rp_data                 (rsp_xbar_mux_001_src_data),                                                            //          .data
		.rp_channel              (rsp_xbar_mux_001_src_channel),                                                         //          .channel
		.rp_startofpacket        (rsp_xbar_mux_001_src_startofpacket),                                                   //          .startofpacket
		.rp_endofpacket          (rsp_xbar_mux_001_src_endofpacket),                                                     //          .endofpacket
		.rp_ready                (rsp_xbar_mux_001_src_ready),                                                           //          .ready
		.av_response             (),                                                                                     // (terminated)
		.av_writeresponserequest (1'b0),                                                                                 // (terminated)
		.av_writeresponsevalid   ()                                                                                      // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (82),
		.PKT_PROTECTION_L          (80),
		.PKT_BEGIN_BURST           (69),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.PKT_BURST_TYPE_H          (66),
		.PKT_BURST_TYPE_L          (65),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_TRANS_EXCLUSIVE       (55),
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_SRC_ID_H              (74),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (78),
		.PKT_DEST_ID_L             (75),
		.PKT_THREAD_ID_H           (79),
		.PKT_THREAD_ID_L           (79),
		.PKT_CACHE_H               (86),
		.PKT_CACHE_L               (83),
		.PKT_DATA_SIDEBAND_H       (68),
		.PKT_DATA_SIDEBAND_L       (68),
		.PKT_QOS_H                 (70),
		.PKT_QOS_L                 (70),
		.PKT_ADDR_SIDEBAND_H       (67),
		.PKT_ADDR_SIDEBAND_L       (67),
		.PKT_RESPONSE_STATUS_H     (88),
		.PKT_RESPONSE_STATUS_L     (87),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (16),
		.AV_BURSTCOUNT_W           (2),
		.SUPPRESS_0_BYTEEN_RSP     (1),
		.ID                        (3),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                                   //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                       // clk_reset.reset
		.av_address              (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_demux_010_src1_valid),                                                                        //        rp.valid
		.rp_data                 (rsp_xbar_demux_010_src1_data),                                                                         //          .data
		.rp_channel              (rsp_xbar_demux_010_src1_channel),                                                                      //          .channel
		.rp_startofpacket        (rsp_xbar_demux_010_src1_startofpacket),                                                                //          .startofpacket
		.rp_endofpacket          (rsp_xbar_demux_010_src1_endofpacket),                                                                  //          .endofpacket
		.rp_ready                (rsp_xbar_demux_010_src1_ready),                                                                        //          .ready
		.av_response             (),                                                                                                     // (terminated)
		.av_writeresponserequest (1'b0),                                                                                                 // (terminated)
		.av_writeresponsevalid   ()                                                                                                      // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (82),
		.PKT_PROTECTION_L          (80),
		.PKT_BEGIN_BURST           (69),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.PKT_BURST_TYPE_H          (66),
		.PKT_BURST_TYPE_L          (65),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_TRANS_EXCLUSIVE       (55),
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_SRC_ID_H              (74),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (78),
		.PKT_DEST_ID_L             (75),
		.PKT_THREAD_ID_H           (79),
		.PKT_THREAD_ID_L           (79),
		.PKT_CACHE_H               (86),
		.PKT_CACHE_L               (83),
		.PKT_DATA_SIDEBAND_H       (68),
		.PKT_DATA_SIDEBAND_L       (68),
		.PKT_QOS_H                 (70),
		.PKT_QOS_L                 (70),
		.PKT_ADDR_SIDEBAND_H       (67),
		.PKT_ADDR_SIDEBAND_L       (67),
		.PKT_RESPONSE_STATUS_H     (88),
		.PKT_RESPONSE_STATUS_L     (87),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (16),
		.AV_BURSTCOUNT_W           (2),
		.SUPPRESS_0_BYTEEN_RSP     (1),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) line_drawer_0_avalon_master_translator_avalon_universal_master_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                      //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                          // clk_reset.reset
		.av_address              (line_drawer_0_avalon_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (line_drawer_0_avalon_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (line_drawer_0_avalon_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (line_drawer_0_avalon_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (line_drawer_0_avalon_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (line_drawer_0_avalon_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (line_drawer_0_avalon_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (line_drawer_0_avalon_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (line_drawer_0_avalon_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (line_drawer_0_avalon_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (line_drawer_0_avalon_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (line_drawer_0_avalon_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (line_drawer_0_avalon_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (line_drawer_0_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (line_drawer_0_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (line_drawer_0_avalon_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_demux_010_src2_valid),                                                           //        rp.valid
		.rp_data                 (rsp_xbar_demux_010_src2_data),                                                            //          .data
		.rp_channel              (rsp_xbar_demux_010_src2_channel),                                                         //          .channel
		.rp_startofpacket        (rsp_xbar_demux_010_src2_startofpacket),                                                   //          .startofpacket
		.rp_endofpacket          (rsp_xbar_demux_010_src2_endofpacket),                                                     //          .endofpacket
		.rp_ready                (rsp_xbar_demux_010_src2_ready),                                                           //          .ready
		.av_response             (),                                                                                        // (terminated)
		.av_writeresponserequest (1'b0),                                                                                    // (terminated)
		.av_writeresponsevalid   ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                                  //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                      //       clk_reset.reset
		.m0_address              (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                              //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                              //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                               //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                                      //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                                        //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                            //                .channel
		.rf_sink_ready           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                               //     (terminated)
		.m0_writeresponserequest (),                                                                                                    //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                 //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                                  //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                      // clk_reset.reset
		.in_data           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                                // (terminated)
		.csr_readdata      (),                                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                // (terminated)
		.almost_full_data  (),                                                                                                    // (terminated)
		.almost_empty_data (),                                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                                // (terminated)
		.out_empty         (),                                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                                // (terminated)
		.out_error         (),                                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                                // (terminated)
		.out_channel       ()                                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                       //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_001_src_ready),                                                               //              cp.ready
		.cp_valid                (cmd_xbar_mux_001_src_valid),                                                               //                .valid
		.cp_data                 (cmd_xbar_mux_001_src_data),                                                                //                .data
		.cp_startofpacket        (cmd_xbar_mux_001_src_startofpacket),                                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_001_src_endofpacket),                                                         //                .endofpacket
		.cp_channel              (cmd_xbar_mux_001_src_channel),                                                             //                .channel
		.rf_sink_ready           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                    //     (terminated)
		.m0_writeresponserequest (),                                                                                         //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                      //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                       //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (74),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (78),
		.PKT_DEST_ID_L             (75),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (82),
		.PKT_PROTECTION_L          (80),
		.PKT_RESPONSE_STATUS_H     (88),
		.PKT_RESPONSE_STATUS_L     (87),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (89),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sdram_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                            //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (sdram_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sdram_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sdram_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_source0_ready),                                                   //              cp.ready
		.cp_valid                (burst_adapter_source0_valid),                                                   //                .valid
		.cp_data                 (burst_adapter_source0_data),                                                    //                .data
		.cp_startofpacket        (burst_adapter_source0_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (burst_adapter_source0_endofpacket),                                             //                .endofpacket
		.cp_channel              (burst_adapter_source0_channel),                                                 //                .channel
		.rf_sink_ready           (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (90),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                            //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.in_data           (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (18),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clocks_sys_clk_clk),                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                          // clk_reset.reset
		.in_data           (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                   // (terminated)
		.csr_read          (1'b0),                                                                    // (terminated)
		.csr_write         (1'b0),                                                                    // (terminated)
		.csr_readdata      (),                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                    // (terminated)
		.almost_full_data  (),                                                                        // (terminated)
		.almost_empty_data (),                                                                        // (terminated)
		.in_startofpacket  (1'b0),                                                                    // (terminated)
		.in_endofpacket    (1'b0),                                                                    // (terminated)
		.out_startofpacket (),                                                                        // (terminated)
		.out_endofpacket   (),                                                                        // (terminated)
		.in_empty          (1'b0),                                                                    // (terminated)
		.out_empty         (),                                                                        // (terminated)
		.in_error          (1'b0),                                                                    // (terminated)
		.out_error         (),                                                                        // (terminated)
		.in_channel        (1'b0),                                                                    // (terminated)
		.out_channel       ()                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) timer_system_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                   //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                       //       clk_reset.reset
		.m0_address              (timer_system_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_system_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_system_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_system_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_system_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_system_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_system_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_system_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_system_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_system_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_system_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_system_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_system_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_system_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_system_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_system_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_003_src_ready),                                                           //              cp.ready
		.cp_valid                (cmd_xbar_mux_003_src_valid),                                                           //                .valid
		.cp_data                 (cmd_xbar_mux_003_src_data),                                                            //                .data
		.cp_startofpacket        (cmd_xbar_mux_003_src_startofpacket),                                                   //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_003_src_endofpacket),                                                     //                .endofpacket
		.cp_channel              (cmd_xbar_mux_003_src_channel),                                                         //                .channel
		.rf_sink_ready           (timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_system_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_system_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_system_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_system_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_system_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_system_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_system_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_system_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timer_system_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_system_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_system_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                //     (terminated)
		.m0_writeresponserequest (),                                                                                     //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                  //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                   //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.in_data           (timer_system_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_system_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_system_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_system_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_system_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_system_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                // (terminated)
		.csr_read          (1'b0),                                                                                 // (terminated)
		.csr_write         (1'b0),                                                                                 // (terminated)
		.csr_readdata      (),                                                                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                 // (terminated)
		.almost_full_data  (),                                                                                     // (terminated)
		.almost_empty_data (),                                                                                     // (terminated)
		.in_empty          (1'b0),                                                                                 // (terminated)
		.out_empty         (),                                                                                     // (terminated)
		.in_error          (1'b0),                                                                                 // (terminated)
		.out_error         (),                                                                                     // (terminated)
		.in_channel        (1'b0),                                                                                 // (terminated)
		.out_channel       ()                                                                                      // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) timer_timestamp_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                      //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                          //       clk_reset.reset
		.m0_address              (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_004_src_ready),                                                              //              cp.ready
		.cp_valid                (cmd_xbar_mux_004_src_valid),                                                              //                .valid
		.cp_data                 (cmd_xbar_mux_004_src_data),                                                               //                .data
		.cp_startofpacket        (cmd_xbar_mux_004_src_startofpacket),                                                      //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_004_src_endofpacket),                                                        //                .endofpacket
		.cp_channel              (cmd_xbar_mux_004_src_channel),                                                            //                .channel
		.rf_sink_ready           (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                   //     (terminated)
		.m0_writeresponserequest (),                                                                                        //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                     //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                          // clk_reset.reset
		.in_data           (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                               //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                   //       clk_reset.reset
		.m0_address              (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_005_src_ready),                                                                       //              cp.ready
		.cp_valid                (cmd_xbar_mux_005_src_valid),                                                                       //                .valid
		.cp_data                 (cmd_xbar_mux_005_src_data),                                                                        //                .data
		.cp_startofpacket        (cmd_xbar_mux_005_src_startofpacket),                                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_005_src_endofpacket),                                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_mux_005_src_channel),                                                                     //                .channel
		.rf_sink_ready           (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                               //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                   // clk_reset.reset
		.in_data           (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                            // (terminated)
		.csr_read          (1'b0),                                                                                             // (terminated)
		.csr_write         (1'b0),                                                                                             // (terminated)
		.csr_readdata      (),                                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                             // (terminated)
		.almost_full_data  (),                                                                                                 // (terminated)
		.almost_empty_data (),                                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                                             // (terminated)
		.out_empty         (),                                                                                                 // (terminated)
		.in_error          (1'b0),                                                                                             // (terminated)
		.out_error         (),                                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                                             // (terminated)
		.out_channel       ()                                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) keys_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                           //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (keys_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (keys_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (keys_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (keys_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (keys_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (keys_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (keys_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (keys_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (keys_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (keys_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (keys_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (keys_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (keys_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (keys_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (keys_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (keys_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src6_ready),                                                //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src6_valid),                                                //                .valid
		.cp_data                 (cmd_xbar_demux_001_src6_data),                                                 //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src6_startofpacket),                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src6_endofpacket),                                          //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src6_channel),                                              //                .channel
		.rf_sink_ready           (keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (keys_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (keys_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (keys_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (keys_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (keys_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (keys_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (keys_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (keys_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (keys_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (keys_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (keys_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (keys_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (keys_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (keys_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (keys_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (keys_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) leds_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                           //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (leds_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (leds_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (leds_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (leds_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (leds_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (leds_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (leds_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (leds_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (leds_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (leds_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (leds_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (leds_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (leds_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (leds_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (leds_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (leds_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src7_ready),                                                //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src7_valid),                                                //                .valid
		.cp_data                 (cmd_xbar_demux_001_src7_data),                                                 //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src7_startofpacket),                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src7_endofpacket),                                          //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src7_channel),                                              //                .channel
		.rf_sink_ready           (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                     //       clk_reset.reset
		.m0_address              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src8_ready),                                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src8_valid),                                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_001_src8_data),                                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src8_startofpacket),                                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src8_endofpacket),                                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src8_channel),                                                                    //                .channel
		.rf_sink_ready           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                     // clk_reset.reset
		.in_data           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                              // (terminated)
		.csr_read          (1'b0),                                                                                               // (terminated)
		.csr_write         (1'b0),                                                                                               // (terminated)
		.csr_readdata      (),                                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                               // (terminated)
		.almost_full_data  (),                                                                                                   // (terminated)
		.almost_empty_data (),                                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                                               // (terminated)
		.out_empty         (),                                                                                                   // (terminated)
		.in_error          (1'b0),                                                                                               // (terminated)
		.out_error         (),                                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                                               // (terminated)
		.out_channel       ()                                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (60),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (65),
		.PKT_SRC_ID_L              (62),
		.PKT_DEST_ID_H             (69),
		.PKT_DEST_ID_L             (66),
		.PKT_BURSTWRAP_H           (52),
		.PKT_BURSTWRAP_L           (50),
		.PKT_BYTE_CNT_H            (49),
		.PKT_BYTE_CNT_L            (47),
		.PKT_PROTECTION_H          (73),
		.PKT_PROTECTION_L          (71),
		.PKT_RESPONSE_STATUS_H     (79),
		.PKT_RESPONSE_STATUS_L     (78),
		.PKT_BURST_SIZE_H          (55),
		.PKT_BURST_SIZE_L          (53),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (80),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                                    //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                        //       clk_reset.reset
		.m0_address              (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_001_source0_ready),                                                                       //              cp.ready
		.cp_valid                (burst_adapter_001_source0_valid),                                                                       //                .valid
		.cp_data                 (burst_adapter_001_source0_data),                                                                        //                .data
		.cp_startofpacket        (burst_adapter_001_source0_startofpacket),                                                               //                .startofpacket
		.cp_endofpacket          (burst_adapter_001_source0_endofpacket),                                                                 //                .endofpacket
		.cp_channel              (burst_adapter_001_source0_channel),                                                                     //                .channel
		.rf_sink_ready           (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                 //     (terminated)
		.m0_writeresponserequest (),                                                                                                      //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                   //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (81),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                                    //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                        // clk_reset.reset
		.in_data           (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                                  // (terminated)
		.csr_readdata      (),                                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                  // (terminated)
		.almost_full_data  (),                                                                                                      // (terminated)
		.almost_empty_data (),                                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                                  // (terminated)
		.out_empty         (),                                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                                  // (terminated)
		.out_error         (),                                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                                  // (terminated)
		.out_channel       ()                                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (74),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (78),
		.PKT_DEST_ID_L             (75),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (82),
		.PKT_PROTECTION_L          (80),
		.PKT_RESPONSE_STATUS_H     (88),
		.PKT_RESPONSE_STATUS_L     (87),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (89),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                                  //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                      //       clk_reset.reset
		.m0_address              (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_002_source0_ready),                                                                     //              cp.ready
		.cp_valid                (burst_adapter_002_source0_valid),                                                                     //                .valid
		.cp_data                 (burst_adapter_002_source0_data),                                                                      //                .data
		.cp_startofpacket        (burst_adapter_002_source0_startofpacket),                                                             //                .startofpacket
		.cp_endofpacket          (burst_adapter_002_source0_endofpacket),                                                               //                .endofpacket
		.cp_channel              (burst_adapter_002_source0_channel),                                                                   //                .channel
		.rf_sink_ready           (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                               //     (terminated)
		.m0_writeresponserequest (),                                                                                                    //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                 //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (90),
		.FIFO_DEPTH          (3),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                                  //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                      // clk_reset.reset
		.in_data           (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                                // (terminated)
		.csr_readdata      (),                                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                // (terminated)
		.almost_full_data  (),                                                                                                    // (terminated)
		.almost_empty_data (),                                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                                // (terminated)
		.out_empty         (),                                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                                // (terminated)
		.out_error         (),                                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                                // (terminated)
		.out_channel       ()                                                                                                     // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (18),
		.FIFO_DEPTH          (3),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clocks_sys_clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                // clk_reset.reset
		.in_data           (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                         // (terminated)
		.csr_read          (1'b0),                                                                                          // (terminated)
		.csr_write         (1'b0),                                                                                          // (terminated)
		.csr_readdata      (),                                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                          // (terminated)
		.almost_full_data  (),                                                                                              // (terminated)
		.almost_empty_data (),                                                                                              // (terminated)
		.in_startofpacket  (1'b0),                                                                                          // (terminated)
		.in_endofpacket    (1'b0),                                                                                          // (terminated)
		.out_startofpacket (),                                                                                              // (terminated)
		.out_endofpacket   (),                                                                                              // (terminated)
		.in_empty          (1'b0),                                                                                          // (terminated)
		.out_empty         (),                                                                                              // (terminated)
		.in_error          (1'b0),                                                                                          // (terminated)
		.out_error         (),                                                                                              // (terminated)
		.in_channel        (1'b0),                                                                                          // (terminated)
		.out_channel       ()                                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                                         //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                             //       clk_reset.reset
		.m0_address              (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src11_ready),                                                                             //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src11_valid),                                                                             //                .valid
		.cp_data                 (cmd_xbar_demux_001_src11_data),                                                                              //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src11_startofpacket),                                                                     //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src11_endofpacket),                                                                       //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src11_channel),                                                                           //                .channel
		.rf_sink_ready           (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                      //     (terminated)
		.m0_writeresponserequest (),                                                                                                           //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                        //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                                         //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                             // clk_reset.reset
		.in_data           (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                                       // (terminated)
		.csr_readdata      (),                                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                       // (terminated)
		.almost_full_data  (),                                                                                                           // (terminated)
		.almost_empty_data (),                                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                                       // (terminated)
		.out_empty         (),                                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                                       // (terminated)
		.out_error         (),                                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                                       // (terminated)
		.out_channel       ()                                                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                                //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                    //       clk_reset.reset
		.m0_address              (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src12_ready),                                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src12_valid),                                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src12_data),                                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src12_startofpacket),                                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src12_endofpacket),                                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src12_channel),                                                                  //                .channel
		.rf_sink_ready           (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                                //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                    // clk_reset.reset
		.in_data           (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                             // (terminated)
		.csr_read          (1'b0),                                                                                              // (terminated)
		.csr_write         (1'b0),                                                                                              // (terminated)
		.csr_readdata      (),                                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                              // (terminated)
		.almost_full_data  (),                                                                                                  // (terminated)
		.almost_empty_data (),                                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                                              // (terminated)
		.out_empty         (),                                                                                                  // (terminated)
		.in_error          (1'b0),                                                                                              // (terminated)
		.out_error         (),                                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                                              // (terminated)
		.out_channel       ()                                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (60),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (65),
		.PKT_SRC_ID_L              (62),
		.PKT_DEST_ID_H             (69),
		.PKT_DEST_ID_L             (66),
		.PKT_BURSTWRAP_H           (52),
		.PKT_BURSTWRAP_L           (50),
		.PKT_BYTE_CNT_H            (49),
		.PKT_BYTE_CNT_L            (47),
		.PKT_PROTECTION_H          (73),
		.PKT_PROTECTION_L          (71),
		.PKT_RESPONSE_STATUS_H     (79),
		.PKT_RESPONSE_STATUS_L     (78),
		.PKT_BURST_SIZE_H          (55),
		.PKT_BURST_SIZE_L          (53),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (80),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) dual_port_ram_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                    //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_003_source0_ready),                                                       //              cp.ready
		.cp_valid                (burst_adapter_003_source0_valid),                                                       //                .valid
		.cp_data                 (burst_adapter_003_source0_data),                                                        //                .data
		.cp_startofpacket        (burst_adapter_003_source0_startofpacket),                                               //                .startofpacket
		.cp_endofpacket          (burst_adapter_003_source0_endofpacket),                                                 //                .endofpacket
		.cp_channel              (burst_adapter_003_source0_channel),                                                     //                .channel
		.rf_sink_ready           (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                 //     (terminated)
		.m0_writeresponserequest (),                                                                                      //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                   //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (81),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                    //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) pi_request_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (pi_request_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pi_request_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pi_request_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pi_request_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pi_request_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pi_request_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pi_request_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pi_request_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pi_request_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pi_request_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pi_request_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pi_request_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pi_request_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pi_request_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pi_request_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pi_request_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src14_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src14_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src14_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src14_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src14_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src14_channel),                                                   //                .channel
		.rf_sink_ready           (pi_request_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pi_request_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pi_request_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pi_request_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pi_request_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pi_request_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pi_request_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pi_request_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pi_request_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pi_request_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pi_request_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pi_request_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pi_request_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pi_request_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pi_request_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pi_request_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pi_request_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (pi_request_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pi_request_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pi_request_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pi_request_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pi_request_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pi_request_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pi_request_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pi_request_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pi_request_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pi_request_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) de2_ack_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                              //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (de2_ack_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (de2_ack_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (de2_ack_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (de2_ack_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (de2_ack_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (de2_ack_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (de2_ack_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (de2_ack_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (de2_ack_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (de2_ack_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (de2_ack_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (de2_ack_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (de2_ack_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (de2_ack_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (de2_ack_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (de2_ack_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src15_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src15_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src15_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src15_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src15_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src15_channel),                                                //                .channel
		.rf_sink_ready           (de2_ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (de2_ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (de2_ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (de2_ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (de2_ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (de2_ack_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (de2_ack_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (de2_ack_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (de2_ack_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (de2_ack_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (de2_ack_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (de2_ack_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (de2_ack_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (de2_ack_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (de2_ack_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (de2_ack_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) de2_ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                              //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (de2_ack_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (de2_ack_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (de2_ack_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (de2_ack_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (de2_ack_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (de2_ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (de2_ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (de2_ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (de2_ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (de2_ack_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	nios_system_addr_router addr_router (
		.sink_ready         (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                                       //       src.ready
		.src_valid          (addr_router_src_valid),                                                                       //          .valid
		.src_data           (addr_router_src_data),                                                                        //          .data
		.src_channel        (addr_router_src_channel),                                                                     //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                               //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                                  //          .endofpacket
	);

	nios_system_addr_router_001 addr_router_001 (
		.sink_ready         (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                            //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                            //          .valid
		.src_data           (addr_router_001_src_data),                                                             //          .data
		.src_channel        (addr_router_001_src_channel),                                                          //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                       //          .endofpacket
	);

	nios_system_addr_router_002 addr_router_002 (
		.sink_ready         (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                       // clk_reset.reset
		.src_ready          (addr_router_002_src_ready),                                                                            //       src.ready
		.src_valid          (addr_router_002_src_valid),                                                                            //          .valid
		.src_data           (addr_router_002_src_data),                                                                             //          .data
		.src_channel        (addr_router_002_src_channel),                                                                          //          .channel
		.src_startofpacket  (addr_router_002_src_startofpacket),                                                                    //          .startofpacket
		.src_endofpacket    (addr_router_002_src_endofpacket)                                                                       //          .endofpacket
	);

	nios_system_addr_router_002 addr_router_003 (
		.sink_ready         (line_drawer_0_avalon_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (line_drawer_0_avalon_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (line_drawer_0_avalon_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (line_drawer_0_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (line_drawer_0_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                          // clk_reset.reset
		.src_ready          (addr_router_003_src_ready),                                                               //       src.ready
		.src_valid          (addr_router_003_src_valid),                                                               //          .valid
		.src_data           (addr_router_003_src_data),                                                                //          .data
		.src_channel        (addr_router_003_src_channel),                                                             //          .channel
		.src_startofpacket  (addr_router_003_src_startofpacket),                                                       //          .startofpacket
		.src_endofpacket    (addr_router_003_src_endofpacket)                                                          //          .endofpacket
	);

	nios_system_id_router id_router (
		.sink_ready         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                                       //       src.ready
		.src_valid          (id_router_src_valid),                                                                       //          .valid
		.src_data           (id_router_src_data),                                                                        //          .data
		.src_channel        (id_router_src_channel),                                                                     //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                               //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                                  //          .endofpacket
	);

	nios_system_id_router id_router_001 (
		.sink_ready         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                             //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                        //       src.ready
		.src_valid          (id_router_001_src_valid),                                                        //          .valid
		.src_data           (id_router_001_src_data),                                                         //          .data
		.src_channel        (id_router_001_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                                   //          .endofpacket
	);

	nios_system_id_router_002 id_router_002 (
		.sink_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                             //       src.ready
		.src_valid          (id_router_002_src_valid),                                             //          .valid
		.src_data           (id_router_002_src_data),                                              //          .data
		.src_channel        (id_router_002_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                        //          .endofpacket
	);

	nios_system_id_router id_router_003 (
		.sink_ready         (timer_system_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_system_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_system_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_system_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_system_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                             // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                    //       src.ready
		.src_valid          (id_router_003_src_valid),                                                    //          .valid
		.src_data           (id_router_003_src_data),                                                     //          .data
		.src_channel        (id_router_003_src_channel),                                                  //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                            //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                               //          .endofpacket
	);

	nios_system_id_router id_router_004 (
		.sink_ready         (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_timestamp_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                       //       src.ready
		.src_valid          (id_router_004_src_valid),                                                       //          .valid
		.src_data           (id_router_004_src_data),                                                        //          .data
		.src_channel        (id_router_004_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                                  //          .endofpacket
	);

	nios_system_id_router id_router_005 (
		.sink_ready         (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                         // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                                                //       src.ready
		.src_valid          (id_router_005_src_valid),                                                                //          .valid
		.src_data           (id_router_005_src_data),                                                                 //          .data
		.src_channel        (id_router_005_src_channel),                                                              //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                                           //          .endofpacket
	);

	nios_system_id_router_006 id_router_006 (
		.sink_ready         (keys_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (keys_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (keys_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (keys_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (keys_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                            //       src.ready
		.src_valid          (id_router_006_src_valid),                                            //          .valid
		.src_data           (id_router_006_src_data),                                             //          .data
		.src_channel        (id_router_006_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                       //          .endofpacket
	);

	nios_system_id_router_006 id_router_007 (
		.sink_ready         (leds_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (leds_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (leds_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (leds_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (leds_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                            //       src.ready
		.src_valid          (id_router_007_src_valid),                                            //          .valid
		.src_data           (id_router_007_src_data),                                             //          .data
		.src_channel        (id_router_007_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                       //          .endofpacket
	);

	nios_system_id_router_006 id_router_008 (
		.sink_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                                                  //       src.ready
		.src_valid          (id_router_008_src_valid),                                                                  //          .valid
		.src_data           (id_router_008_src_data),                                                                   //          .data
		.src_channel        (id_router_008_src_channel),                                                                //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                                             //          .endofpacket
	);

	nios_system_id_router_009 id_router_009 (
		.sink_ready         (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.src_ready          (id_router_009_src_ready),                                                                     //       src.ready
		.src_valid          (id_router_009_src_valid),                                                                     //          .valid
		.src_data           (id_router_009_src_data),                                                                      //          .data
		.src_channel        (id_router_009_src_channel),                                                                   //          .channel
		.src_startofpacket  (id_router_009_src_startofpacket),                                                             //          .startofpacket
		.src_endofpacket    (id_router_009_src_endofpacket)                                                                //          .endofpacket
	);

	nios_system_id_router_010 id_router_010 (
		.sink_ready         (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.src_ready          (id_router_010_src_ready),                                                                   //       src.ready
		.src_valid          (id_router_010_src_valid),                                                                   //          .valid
		.src_data           (id_router_010_src_data),                                                                    //          .data
		.src_channel        (id_router_010_src_channel),                                                                 //          .channel
		.src_startofpacket  (id_router_010_src_startofpacket),                                                           //          .startofpacket
		.src_endofpacket    (id_router_010_src_endofpacket)                                                              //          .endofpacket
	);

	nios_system_id_router_006 id_router_011 (
		.sink_ready         (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                   // clk_reset.reset
		.src_ready          (id_router_011_src_ready),                                                                          //       src.ready
		.src_valid          (id_router_011_src_valid),                                                                          //          .valid
		.src_data           (id_router_011_src_data),                                                                           //          .data
		.src_channel        (id_router_011_src_channel),                                                                        //          .channel
		.src_startofpacket  (id_router_011_src_startofpacket),                                                                  //          .startofpacket
		.src_endofpacket    (id_router_011_src_endofpacket)                                                                     //          .endofpacket
	);

	nios_system_id_router_006 id_router_012 (
		.sink_ready         (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (line_drawer_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                          // clk_reset.reset
		.src_ready          (id_router_012_src_ready),                                                                 //       src.ready
		.src_valid          (id_router_012_src_valid),                                                                 //          .valid
		.src_data           (id_router_012_src_data),                                                                  //          .data
		.src_channel        (id_router_012_src_channel),                                                               //          .channel
		.src_startofpacket  (id_router_012_src_startofpacket),                                                         //          .startofpacket
		.src_endofpacket    (id_router_012_src_endofpacket)                                                            //          .endofpacket
	);

	nios_system_id_router_009 id_router_013 (
		.sink_ready         (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (dual_port_ram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (id_router_013_src_ready),                                                     //       src.ready
		.src_valid          (id_router_013_src_valid),                                                     //          .valid
		.src_data           (id_router_013_src_data),                                                      //          .data
		.src_channel        (id_router_013_src_channel),                                                   //          .channel
		.src_startofpacket  (id_router_013_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (id_router_013_src_endofpacket)                                                //          .endofpacket
	);

	nios_system_id_router_006 id_router_014 (
		.sink_ready         (pi_request_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pi_request_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pi_request_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pi_request_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pi_request_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_014_src_ready),                                                  //       src.ready
		.src_valid          (id_router_014_src_valid),                                                  //          .valid
		.src_data           (id_router_014_src_data),                                                   //          .data
		.src_channel        (id_router_014_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_014_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_014_src_endofpacket)                                             //          .endofpacket
	);

	nios_system_id_router_006 id_router_015 (
		.sink_ready         (de2_ack_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (de2_ack_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (de2_ack_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (de2_ack_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (de2_ack_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_015_src_ready),                                               //       src.ready
		.src_valid          (id_router_015_src_valid),                                               //          .valid
		.src_data           (id_router_015_src_data),                                                //          .data
		.src_channel        (id_router_015_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_015_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_015_src_endofpacket)                                          //          .endofpacket
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (69),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.PKT_BURST_TYPE_H          (66),
		.PKT_BURST_TYPE_L          (65),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (16),
		.OUT_BYTE_CNT_H            (57),
		.OUT_BURSTWRAP_H           (61),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (3),
		.BURSTWRAP_CONST_VALUE     (3)
	) burst_adapter (
		.clk                   (clocks_sys_clk_clk),                  //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (cmd_xbar_mux_002_src_valid),          //     sink0.valid
		.sink0_data            (cmd_xbar_mux_002_src_data),           //          .data
		.sink0_channel         (cmd_xbar_mux_002_src_channel),        //          .channel
		.sink0_startofpacket   (cmd_xbar_mux_002_src_startofpacket),  //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_mux_002_src_endofpacket),    //          .endofpacket
		.sink0_ready           (cmd_xbar_mux_002_src_ready),          //          .ready
		.source0_valid         (burst_adapter_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_source0_data),          //          .data
		.source0_channel       (burst_adapter_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (60),
		.PKT_BYTE_CNT_H            (49),
		.PKT_BYTE_CNT_L            (47),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURST_SIZE_H          (55),
		.PKT_BURST_SIZE_L          (53),
		.PKT_BURST_TYPE_H          (57),
		.PKT_BURST_TYPE_L          (56),
		.PKT_BURSTWRAP_H           (52),
		.PKT_BURSTWRAP_L           (50),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (80),
		.ST_CHANNEL_W              (16),
		.OUT_BYTE_CNT_H            (47),
		.OUT_BURSTWRAP_H           (52),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_001 (
		.clk                   (clocks_sys_clk_clk),                      //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (width_adapter_002_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_002_src_data),              //          .data
		.sink0_channel         (width_adapter_002_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_002_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_002_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_002_src_ready),             //          .ready
		.source0_valid         (burst_adapter_001_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_001_source0_data),          //          .data
		.source0_channel       (burst_adapter_001_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_001_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_001_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_001_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (69),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.PKT_BURST_TYPE_H          (66),
		.PKT_BURST_TYPE_L          (65),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (16),
		.OUT_BYTE_CNT_H            (57),
		.OUT_BURSTWRAP_H           (61),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_002 (
		.clk                   (clocks_sys_clk_clk),                      //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (cmd_xbar_mux_010_src_valid),              //     sink0.valid
		.sink0_data            (cmd_xbar_mux_010_src_data),               //          .data
		.sink0_channel         (cmd_xbar_mux_010_src_channel),            //          .channel
		.sink0_startofpacket   (cmd_xbar_mux_010_src_startofpacket),      //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_mux_010_src_endofpacket),        //          .endofpacket
		.sink0_ready           (cmd_xbar_mux_010_src_ready),              //          .ready
		.source0_valid         (burst_adapter_002_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_002_source0_data),          //          .data
		.source0_channel       (burst_adapter_002_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_002_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_002_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_002_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (60),
		.PKT_BYTE_CNT_H            (49),
		.PKT_BYTE_CNT_L            (47),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURST_SIZE_H          (55),
		.PKT_BURST_SIZE_L          (53),
		.PKT_BURST_TYPE_H          (57),
		.PKT_BURST_TYPE_L          (56),
		.PKT_BURSTWRAP_H           (52),
		.PKT_BURSTWRAP_L           (50),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (80),
		.ST_CHANNEL_W              (16),
		.OUT_BYTE_CNT_H            (47),
		.OUT_BURSTWRAP_H           (52),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_003 (
		.clk                   (clocks_sys_clk_clk),                      //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (width_adapter_004_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_004_src_data),              //          .data
		.sink0_channel         (width_adapter_004_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_004_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_004_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_004_src_ready),             //          .ready
		.source0_valid         (burst_adapter_003_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_003_source0_data),          //          .data
		.source0_channel       (burst_adapter_003_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_003_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_003_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_003_source0_ready)          //          .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (1)
	) rst_controller (
		.reset_in0  (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in0.reset
		.reset_in1  (~reset_reset_n),                             // reset_in1.reset
		.clk        (clocks_sys_clk_clk),                         //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),             // reset_out.reset
		.reset_req  (rst_controller_reset_out_reset_req),         //          .reset_req
		.reset_in2  (1'b0),                                       // (terminated)
		.reset_in3  (1'b0),                                       // (terminated)
		.reset_in4  (1'b0),                                       // (terminated)
		.reset_in5  (1'b0),                                       // (terminated)
		.reset_in6  (1'b0),                                       // (terminated)
		.reset_in7  (1'b0),                                       // (terminated)
		.reset_in8  (1'b0),                                       // (terminated)
		.reset_in9  (1'b0),                                       // (terminated)
		.reset_in10 (1'b0),                                       // (terminated)
		.reset_in11 (1'b0),                                       // (terminated)
		.reset_in12 (1'b0),                                       // (terminated)
		.reset_in13 (1'b0),                                       // (terminated)
		.reset_in14 (1'b0),                                       // (terminated)
		.reset_in15 (1'b0)                                        // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_001 (
		.reset_in0  (~reset_reset_n),                             // reset_in0.reset
		.reset_in1  (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (clk_clk),                                    //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset),         // reset_out.reset
		.reset_req  (),                                           // (terminated)
		.reset_in2  (1'b0),                                       // (terminated)
		.reset_in3  (1'b0),                                       // (terminated)
		.reset_in4  (1'b0),                                       // (terminated)
		.reset_in5  (1'b0),                                       // (terminated)
		.reset_in6  (1'b0),                                       // (terminated)
		.reset_in7  (1'b0),                                       // (terminated)
		.reset_in8  (1'b0),                                       // (terminated)
		.reset_in9  (1'b0),                                       // (terminated)
		.reset_in10 (1'b0),                                       // (terminated)
		.reset_in11 (1'b0),                                       // (terminated)
		.reset_in12 (1'b0),                                       // (terminated)
		.reset_in13 (1'b0),                                       // (terminated)
		.reset_in14 (1'b0),                                       // (terminated)
		.reset_in15 (1'b0)                                        // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_002 (
		.reset_in0  (~reset_reset_n),                             // reset_in0.reset
		.reset_in1  (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (clocks_vga_clk_clk),                         //       clk.clk
		.reset_out  (rst_controller_002_reset_out_reset),         // reset_out.reset
		.reset_req  (),                                           // (terminated)
		.reset_in2  (1'b0),                                       // (terminated)
		.reset_in3  (1'b0),                                       // (terminated)
		.reset_in4  (1'b0),                                       // (terminated)
		.reset_in5  (1'b0),                                       // (terminated)
		.reset_in6  (1'b0),                                       // (terminated)
		.reset_in7  (1'b0),                                       // (terminated)
		.reset_in8  (1'b0),                                       // (terminated)
		.reset_in9  (1'b0),                                       // (terminated)
		.reset_in10 (1'b0),                                       // (terminated)
		.reset_in11 (1'b0),                                       // (terminated)
		.reset_in12 (1'b0),                                       // (terminated)
		.reset_in13 (1'b0),                                       // (terminated)
		.reset_in14 (1'b0),                                       // (terminated)
		.reset_in15 (1'b0)                                        // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (3),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (1)
	) rst_controller_003 (
		.reset_in0  (~reset_reset_n),                             // reset_in0.reset
		.reset_in1  (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2  (rst_controller_004_reset_out_reset),         // reset_in2.reset
		.clk        (clk_pi_clk),                                 //       clk.clk
		.reset_out  (rst_controller_003_reset_out_reset),         // reset_out.reset
		.reset_req  (rst_controller_003_reset_out_reset_req),     //          .reset_req
		.reset_in3  (1'b0),                                       // (terminated)
		.reset_in4  (1'b0),                                       // (terminated)
		.reset_in5  (1'b0),                                       // (terminated)
		.reset_in6  (1'b0),                                       // (terminated)
		.reset_in7  (1'b0),                                       // (terminated)
		.reset_in8  (1'b0),                                       // (terminated)
		.reset_in9  (1'b0),                                       // (terminated)
		.reset_in10 (1'b0),                                       // (terminated)
		.reset_in11 (1'b0),                                       // (terminated)
		.reset_in12 (1'b0),                                       // (terminated)
		.reset_in13 (1'b0),                                       // (terminated)
		.reset_in14 (1'b0),                                       // (terminated)
		.reset_in15 (1'b0)                                        // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("none"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_004 (
		.reset_in0  (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in0.reset
		.reset_in1  (~reset_reset_n),                             // reset_in1.reset
		.clk        (),                                           //       clk.clk
		.reset_out  (rst_controller_004_reset_out_reset),         // reset_out.reset
		.reset_req  (),                                           // (terminated)
		.reset_in2  (1'b0),                                       // (terminated)
		.reset_in3  (1'b0),                                       // (terminated)
		.reset_in4  (1'b0),                                       // (terminated)
		.reset_in5  (1'b0),                                       // (terminated)
		.reset_in6  (1'b0),                                       // (terminated)
		.reset_in7  (1'b0),                                       // (terminated)
		.reset_in8  (1'b0),                                       // (terminated)
		.reset_in9  (1'b0),                                       // (terminated)
		.reset_in10 (1'b0),                                       // (terminated)
		.reset_in11 (1'b0),                                       // (terminated)
		.reset_in12 (1'b0),                                       // (terminated)
		.reset_in13 (1'b0),                                       // (terminated)
		.reset_in14 (1'b0),                                       // (terminated)
		.reset_in15 (1'b0)                                        // (terminated)
	);

	nios_system_cmd_xbar_demux cmd_xbar_demux (
		.clk                (clocks_sys_clk_clk),                //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_src_ready),             //      sink.ready
		.sink_channel       (addr_router_src_channel),           //          .channel
		.sink_data          (addr_router_src_data),              //          .data
		.sink_startofpacket (addr_router_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket),   //          .endofpacket
		.src2_ready         (cmd_xbar_demux_src2_ready),         //      src2.ready
		.src2_valid         (cmd_xbar_demux_src2_valid),         //          .valid
		.src2_data          (cmd_xbar_demux_src2_data),          //          .data
		.src2_channel       (cmd_xbar_demux_src2_channel),       //          .channel
		.src2_startofpacket (cmd_xbar_demux_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_src2_endofpacket),   //          .endofpacket
		.src3_ready         (cmd_xbar_demux_src3_ready),         //      src3.ready
		.src3_valid         (cmd_xbar_demux_src3_valid),         //          .valid
		.src3_data          (cmd_xbar_demux_src3_data),          //          .data
		.src3_channel       (cmd_xbar_demux_src3_channel),       //          .channel
		.src3_startofpacket (cmd_xbar_demux_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_src3_endofpacket),   //          .endofpacket
		.src4_ready         (cmd_xbar_demux_src4_ready),         //      src4.ready
		.src4_valid         (cmd_xbar_demux_src4_valid),         //          .valid
		.src4_data          (cmd_xbar_demux_src4_data),          //          .data
		.src4_channel       (cmd_xbar_demux_src4_channel),       //          .channel
		.src4_startofpacket (cmd_xbar_demux_src4_startofpacket), //          .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_src4_endofpacket),   //          .endofpacket
		.src5_ready         (cmd_xbar_demux_src5_ready),         //      src5.ready
		.src5_valid         (cmd_xbar_demux_src5_valid),         //          .valid
		.src5_data          (cmd_xbar_demux_src5_data),          //          .data
		.src5_channel       (cmd_xbar_demux_src5_channel),       //          .channel
		.src5_startofpacket (cmd_xbar_demux_src5_startofpacket), //          .startofpacket
		.src5_endofpacket   (cmd_xbar_demux_src5_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                 (clocks_sys_clk_clk),                     //       clk.clk
		.reset               (rst_controller_reset_out_reset),         // clk_reset.reset
		.sink_ready          (addr_router_001_src_ready),              //      sink.ready
		.sink_channel        (addr_router_001_src_channel),            //          .channel
		.sink_data           (addr_router_001_src_data),               //          .data
		.sink_startofpacket  (addr_router_001_src_startofpacket),      //          .startofpacket
		.sink_endofpacket    (addr_router_001_src_endofpacket),        //          .endofpacket
		.sink_valid          (addr_router_001_src_valid),              //          .valid
		.src0_ready          (cmd_xbar_demux_001_src0_ready),          //      src0.ready
		.src0_valid          (cmd_xbar_demux_001_src0_valid),          //          .valid
		.src0_data           (cmd_xbar_demux_001_src0_data),           //          .data
		.src0_channel        (cmd_xbar_demux_001_src0_channel),        //          .channel
		.src0_startofpacket  (cmd_xbar_demux_001_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_001_src0_endofpacket),    //          .endofpacket
		.src1_ready          (cmd_xbar_demux_001_src1_ready),          //      src1.ready
		.src1_valid          (cmd_xbar_demux_001_src1_valid),          //          .valid
		.src1_data           (cmd_xbar_demux_001_src1_data),           //          .data
		.src1_channel        (cmd_xbar_demux_001_src1_channel),        //          .channel
		.src1_startofpacket  (cmd_xbar_demux_001_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_001_src1_endofpacket),    //          .endofpacket
		.src2_ready          (cmd_xbar_demux_001_src2_ready),          //      src2.ready
		.src2_valid          (cmd_xbar_demux_001_src2_valid),          //          .valid
		.src2_data           (cmd_xbar_demux_001_src2_data),           //          .data
		.src2_channel        (cmd_xbar_demux_001_src2_channel),        //          .channel
		.src2_startofpacket  (cmd_xbar_demux_001_src2_startofpacket),  //          .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_001_src2_endofpacket),    //          .endofpacket
		.src3_ready          (cmd_xbar_demux_001_src3_ready),          //      src3.ready
		.src3_valid          (cmd_xbar_demux_001_src3_valid),          //          .valid
		.src3_data           (cmd_xbar_demux_001_src3_data),           //          .data
		.src3_channel        (cmd_xbar_demux_001_src3_channel),        //          .channel
		.src3_startofpacket  (cmd_xbar_demux_001_src3_startofpacket),  //          .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_001_src3_endofpacket),    //          .endofpacket
		.src4_ready          (cmd_xbar_demux_001_src4_ready),          //      src4.ready
		.src4_valid          (cmd_xbar_demux_001_src4_valid),          //          .valid
		.src4_data           (cmd_xbar_demux_001_src4_data),           //          .data
		.src4_channel        (cmd_xbar_demux_001_src4_channel),        //          .channel
		.src4_startofpacket  (cmd_xbar_demux_001_src4_startofpacket),  //          .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_001_src4_endofpacket),    //          .endofpacket
		.src5_ready          (cmd_xbar_demux_001_src5_ready),          //      src5.ready
		.src5_valid          (cmd_xbar_demux_001_src5_valid),          //          .valid
		.src5_data           (cmd_xbar_demux_001_src5_data),           //          .data
		.src5_channel        (cmd_xbar_demux_001_src5_channel),        //          .channel
		.src5_startofpacket  (cmd_xbar_demux_001_src5_startofpacket),  //          .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_001_src5_endofpacket),    //          .endofpacket
		.src6_ready          (cmd_xbar_demux_001_src6_ready),          //      src6.ready
		.src6_valid          (cmd_xbar_demux_001_src6_valid),          //          .valid
		.src6_data           (cmd_xbar_demux_001_src6_data),           //          .data
		.src6_channel        (cmd_xbar_demux_001_src6_channel),        //          .channel
		.src6_startofpacket  (cmd_xbar_demux_001_src6_startofpacket),  //          .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_001_src6_endofpacket),    //          .endofpacket
		.src7_ready          (cmd_xbar_demux_001_src7_ready),          //      src7.ready
		.src7_valid          (cmd_xbar_demux_001_src7_valid),          //          .valid
		.src7_data           (cmd_xbar_demux_001_src7_data),           //          .data
		.src7_channel        (cmd_xbar_demux_001_src7_channel),        //          .channel
		.src7_startofpacket  (cmd_xbar_demux_001_src7_startofpacket),  //          .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_001_src7_endofpacket),    //          .endofpacket
		.src8_ready          (cmd_xbar_demux_001_src8_ready),          //      src8.ready
		.src8_valid          (cmd_xbar_demux_001_src8_valid),          //          .valid
		.src8_data           (cmd_xbar_demux_001_src8_data),           //          .data
		.src8_channel        (cmd_xbar_demux_001_src8_channel),        //          .channel
		.src8_startofpacket  (cmd_xbar_demux_001_src8_startofpacket),  //          .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_001_src8_endofpacket),    //          .endofpacket
		.src9_ready          (cmd_xbar_demux_001_src9_ready),          //      src9.ready
		.src9_valid          (cmd_xbar_demux_001_src9_valid),          //          .valid
		.src9_data           (cmd_xbar_demux_001_src9_data),           //          .data
		.src9_channel        (cmd_xbar_demux_001_src9_channel),        //          .channel
		.src9_startofpacket  (cmd_xbar_demux_001_src9_startofpacket),  //          .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_001_src9_endofpacket),    //          .endofpacket
		.src10_ready         (cmd_xbar_demux_001_src10_ready),         //     src10.ready
		.src10_valid         (cmd_xbar_demux_001_src10_valid),         //          .valid
		.src10_data          (cmd_xbar_demux_001_src10_data),          //          .data
		.src10_channel       (cmd_xbar_demux_001_src10_channel),       //          .channel
		.src10_startofpacket (cmd_xbar_demux_001_src10_startofpacket), //          .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_001_src10_endofpacket),   //          .endofpacket
		.src11_ready         (cmd_xbar_demux_001_src11_ready),         //     src11.ready
		.src11_valid         (cmd_xbar_demux_001_src11_valid),         //          .valid
		.src11_data          (cmd_xbar_demux_001_src11_data),          //          .data
		.src11_channel       (cmd_xbar_demux_001_src11_channel),       //          .channel
		.src11_startofpacket (cmd_xbar_demux_001_src11_startofpacket), //          .startofpacket
		.src11_endofpacket   (cmd_xbar_demux_001_src11_endofpacket),   //          .endofpacket
		.src12_ready         (cmd_xbar_demux_001_src12_ready),         //     src12.ready
		.src12_valid         (cmd_xbar_demux_001_src12_valid),         //          .valid
		.src12_data          (cmd_xbar_demux_001_src12_data),          //          .data
		.src12_channel       (cmd_xbar_demux_001_src12_channel),       //          .channel
		.src12_startofpacket (cmd_xbar_demux_001_src12_startofpacket), //          .startofpacket
		.src12_endofpacket   (cmd_xbar_demux_001_src12_endofpacket),   //          .endofpacket
		.src13_ready         (cmd_xbar_demux_001_src13_ready),         //     src13.ready
		.src13_valid         (cmd_xbar_demux_001_src13_valid),         //          .valid
		.src13_data          (cmd_xbar_demux_001_src13_data),          //          .data
		.src13_channel       (cmd_xbar_demux_001_src13_channel),       //          .channel
		.src13_startofpacket (cmd_xbar_demux_001_src13_startofpacket), //          .startofpacket
		.src13_endofpacket   (cmd_xbar_demux_001_src13_endofpacket),   //          .endofpacket
		.src14_ready         (cmd_xbar_demux_001_src14_ready),         //     src14.ready
		.src14_valid         (cmd_xbar_demux_001_src14_valid),         //          .valid
		.src14_data          (cmd_xbar_demux_001_src14_data),          //          .data
		.src14_channel       (cmd_xbar_demux_001_src14_channel),       //          .channel
		.src14_startofpacket (cmd_xbar_demux_001_src14_startofpacket), //          .startofpacket
		.src14_endofpacket   (cmd_xbar_demux_001_src14_endofpacket),   //          .endofpacket
		.src15_ready         (cmd_xbar_demux_001_src15_ready),         //     src15.ready
		.src15_valid         (cmd_xbar_demux_001_src15_valid),         //          .valid
		.src15_data          (cmd_xbar_demux_001_src15_data),          //          .data
		.src15_channel       (cmd_xbar_demux_001_src15_channel),       //          .channel
		.src15_startofpacket (cmd_xbar_demux_001_src15_startofpacket), //          .startofpacket
		.src15_endofpacket   (cmd_xbar_demux_001_src15_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_demux_002 cmd_xbar_demux_002 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_002_src_ready),             //      sink.ready
		.sink_channel       (addr_router_002_src_channel),           //          .channel
		.sink_data          (addr_router_002_src_data),              //          .data
		.sink_startofpacket (addr_router_002_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_002_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_002_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_demux_002 cmd_xbar_demux_003 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_003_src_ready),             //      sink.ready
		.sink_channel       (addr_router_003_src_channel),           //          .channel
		.sink_data          (addr_router_003_src_data),              //          .data
		.sink_startofpacket (addr_router_003_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_003_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_003_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (clocks_sys_clk_clk),                    //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux cmd_xbar_mux_001 (
		.clk                 (clocks_sys_clk_clk),                    //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux_002 cmd_xbar_mux_002 (
		.clk                 (clocks_sys_clk_clk),                  //       clk.clk
		.reset               (rst_controller_reset_out_reset),      // clk_reset.reset
		.src_ready           (cmd_xbar_mux_002_src_ready),          //       src.ready
		.src_valid           (cmd_xbar_mux_002_src_valid),          //          .valid
		.src_data            (cmd_xbar_mux_002_src_data),           //          .data
		.src_channel         (cmd_xbar_mux_002_src_channel),        //          .channel
		.src_startofpacket   (cmd_xbar_mux_002_src_startofpacket),  //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_002_src_endofpacket),    //          .endofpacket
		.sink0_ready         (width_adapter_src_ready),             //     sink0.ready
		.sink0_valid         (width_adapter_src_valid),             //          .valid
		.sink0_channel       (width_adapter_src_channel),           //          .channel
		.sink0_data          (width_adapter_src_data),              //          .data
		.sink0_startofpacket (width_adapter_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (width_adapter_src_endofpacket),       //          .endofpacket
		.sink1_ready         (width_adapter_001_src_ready),         //     sink1.ready
		.sink1_valid         (width_adapter_001_src_valid),         //          .valid
		.sink1_channel       (width_adapter_001_src_channel),       //          .channel
		.sink1_data          (width_adapter_001_src_data),          //          .data
		.sink1_startofpacket (width_adapter_001_src_startofpacket), //          .startofpacket
		.sink1_endofpacket   (width_adapter_001_src_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux cmd_xbar_mux_003 (
		.clk                 (clocks_sys_clk_clk),                    //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_003_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_003_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_003_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_003_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_003_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_003_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src3_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src3_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src3_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src3_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src3_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src3_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src3_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src3_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src3_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src3_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src3_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src3_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux cmd_xbar_mux_004 (
		.clk                 (clocks_sys_clk_clk),                    //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_004_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_004_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_004_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_004_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_004_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_004_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src4_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src4_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src4_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src4_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src4_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src4_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src4_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src4_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src4_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src4_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src4_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src4_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux cmd_xbar_mux_005 (
		.clk                 (clocks_sys_clk_clk),                    //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_005_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_005_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_005_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_005_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_005_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_005_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src5_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src5_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src5_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src5_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src5_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src5_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src5_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src5_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src5_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src5_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src5_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src5_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux_010 cmd_xbar_mux_010 (
		.clk                 (clocks_sys_clk_clk),                    //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_010_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_010_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_010_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_010_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_010_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_010_src_endofpacket),      //          .endofpacket
		.sink0_ready         (width_adapter_003_src_ready),           //     sink0.ready
		.sink0_valid         (width_adapter_003_src_valid),           //          .valid
		.sink0_channel       (width_adapter_003_src_channel),         //          .channel
		.sink0_data          (width_adapter_003_src_data),            //          .data
		.sink0_startofpacket (width_adapter_003_src_startofpacket),   //          .startofpacket
		.sink0_endofpacket   (width_adapter_003_src_endofpacket),     //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_002_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_003_src0_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_003_src0_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_003_src0_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_003_src0_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux rsp_xbar_demux (
		.clk                (clocks_sys_clk_clk),                //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_002 rsp_xbar_demux_002 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_002_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_002_src1_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux rsp_xbar_demux_003 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_003_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_003_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_003_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_003_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_003_src1_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux rsp_xbar_demux_004 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_004_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_004_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_004_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_004_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_004_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_004_src1_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux rsp_xbar_demux_005 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_005_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_005_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_005_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_005_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_005_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_005_src1_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_006 rsp_xbar_demux_006 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_006 rsp_xbar_demux_007 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_006 rsp_xbar_demux_008 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_009 rsp_xbar_demux_009 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_009_src_ready),               //      sink.ready
		.sink_channel       (id_router_009_src_channel),             //          .channel
		.sink_data          (id_router_009_src_data),                //          .data
		.sink_startofpacket (id_router_009_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_009_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_009_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_009_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_010 rsp_xbar_demux_010 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_010_src_ready),               //      sink.ready
		.sink_channel       (id_router_010_src_channel),             //          .channel
		.sink_data          (id_router_010_src_data),                //          .data
		.sink_startofpacket (id_router_010_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_010_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_010_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_010_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_010_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_010_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_010_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_010_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_010_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_010_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_010_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_010_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_010_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_010_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_010_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_010_src2_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_006 rsp_xbar_demux_011 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_011_src_ready),               //      sink.ready
		.sink_channel       (id_router_011_src_channel),             //          .channel
		.sink_data          (id_router_011_src_data),                //          .data
		.sink_startofpacket (id_router_011_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_011_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_011_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_011_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_011_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_006 rsp_xbar_demux_012 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_012_src_ready),               //      sink.ready
		.sink_channel       (id_router_012_src_channel),             //          .channel
		.sink_data          (id_router_012_src_data),                //          .data
		.sink_startofpacket (id_router_012_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_012_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_012_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_012_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_012_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_009 rsp_xbar_demux_013 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_013_src_ready),               //      sink.ready
		.sink_channel       (id_router_013_src_channel),             //          .channel
		.sink_data          (id_router_013_src_data),                //          .data
		.sink_startofpacket (id_router_013_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_013_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_013_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_013_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_013_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_006 rsp_xbar_demux_014 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_014_src_ready),               //      sink.ready
		.sink_channel       (id_router_014_src_channel),             //          .channel
		.sink_data          (id_router_014_src_data),                //          .data
		.sink_startofpacket (id_router_014_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_014_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_014_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_014_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_014_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_006 rsp_xbar_demux_015 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_015_src_ready),               //      sink.ready
		.sink_channel       (id_router_015_src_channel),             //          .channel
		.sink_data          (id_router_015_src_data),                //          .data
		.sink_startofpacket (id_router_015_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_015_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_015_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_015_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_015_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (clocks_sys_clk_clk),                    //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (width_adapter_005_src_ready),           //     sink2.ready
		.sink2_valid         (width_adapter_005_src_valid),           //          .valid
		.sink2_channel       (width_adapter_005_src_channel),         //          .channel
		.sink2_data          (width_adapter_005_src_data),            //          .data
		.sink2_startofpacket (width_adapter_005_src_startofpacket),   //          .startofpacket
		.sink2_endofpacket   (width_adapter_005_src_endofpacket),     //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready         (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket   (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink5_ready         (rsp_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                  (clocks_sys_clk_clk),                    //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready            (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel        (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data           (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket  (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready          (width_adapter_006_src_ready),           //     sink2.ready
		.sink2_valid          (width_adapter_006_src_valid),           //          .valid
		.sink2_channel        (width_adapter_006_src_channel),         //          .channel
		.sink2_data           (width_adapter_006_src_data),            //          .data
		.sink2_startofpacket  (width_adapter_006_src_startofpacket),   //          .startofpacket
		.sink2_endofpacket    (width_adapter_006_src_endofpacket),     //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_003_src1_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_003_src1_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_003_src1_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_003_src1_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_003_src1_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_004_src1_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_004_src1_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_004_src1_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_004_src1_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_004_src1_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_004_src1_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_005_src1_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_005_src1_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_005_src1_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_005_src1_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_005_src1_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_005_src1_endofpacket),   //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_006_src0_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_006_src0_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_006_src0_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_006_src0_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_007_src0_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_007_src0_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_007_src0_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_007_src0_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_008_src0_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_008_src0_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_008_src0_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_008_src0_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.sink9_ready          (width_adapter_007_src_ready),           //     sink9.ready
		.sink9_valid          (width_adapter_007_src_valid),           //          .valid
		.sink9_channel        (width_adapter_007_src_channel),         //          .channel
		.sink9_data           (width_adapter_007_src_data),            //          .data
		.sink9_startofpacket  (width_adapter_007_src_startofpacket),   //          .startofpacket
		.sink9_endofpacket    (width_adapter_007_src_endofpacket),     //          .endofpacket
		.sink10_ready         (width_adapter_008_src_ready),           //    sink10.ready
		.sink10_valid         (width_adapter_008_src_valid),           //          .valid
		.sink10_channel       (width_adapter_008_src_channel),         //          .channel
		.sink10_data          (width_adapter_008_src_data),            //          .data
		.sink10_startofpacket (width_adapter_008_src_startofpacket),   //          .startofpacket
		.sink10_endofpacket   (width_adapter_008_src_endofpacket),     //          .endofpacket
		.sink11_ready         (rsp_xbar_demux_011_src0_ready),         //    sink11.ready
		.sink11_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.sink11_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.sink11_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.sink11_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.sink11_endofpacket   (rsp_xbar_demux_011_src0_endofpacket),   //          .endofpacket
		.sink12_ready         (rsp_xbar_demux_012_src0_ready),         //    sink12.ready
		.sink12_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.sink12_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.sink12_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.sink12_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.sink12_endofpacket   (rsp_xbar_demux_012_src0_endofpacket),   //          .endofpacket
		.sink13_ready         (width_adapter_009_src_ready),           //    sink13.ready
		.sink13_valid         (width_adapter_009_src_valid),           //          .valid
		.sink13_channel       (width_adapter_009_src_channel),         //          .channel
		.sink13_data          (width_adapter_009_src_data),            //          .data
		.sink13_startofpacket (width_adapter_009_src_startofpacket),   //          .startofpacket
		.sink13_endofpacket   (width_adapter_009_src_endofpacket),     //          .endofpacket
		.sink14_ready         (rsp_xbar_demux_014_src0_ready),         //    sink14.ready
		.sink14_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.sink14_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.sink14_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.sink14_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.sink14_endofpacket   (rsp_xbar_demux_014_src0_endofpacket),   //          .endofpacket
		.sink15_ready         (rsp_xbar_demux_015_src0_ready),         //    sink15.ready
		.sink15_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.sink15_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.sink15_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.sink15_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.sink15_endofpacket   (rsp_xbar_demux_015_src0_endofpacket)    //          .endofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (106),
		.IN_PKT_RESPONSE_STATUS_L      (105),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (107),
		.OUT_PKT_ADDR_H                (49),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (58),
		.OUT_PKT_BYTE_CNT_L            (56),
		.OUT_PKT_TRANS_COMPRESSED_READ (50),
		.OUT_PKT_BURST_SIZE_H          (64),
		.OUT_PKT_BURST_SIZE_L          (62),
		.OUT_PKT_RESPONSE_STATUS_H     (88),
		.OUT_PKT_RESPONSE_STATUS_L     (87),
		.OUT_PKT_TRANS_EXCLUSIVE       (55),
		.OUT_PKT_BURST_TYPE_H          (66),
		.OUT_PKT_BURST_TYPE_L          (65),
		.OUT_ST_DATA_W                 (89),
		.ST_CHANNEL_W                  (16),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter (
		.clk                  (clocks_sys_clk_clk),                //       clk.clk
		.reset                (rst_controller_reset_out_reset),    // clk_reset.reset
		.in_valid             (cmd_xbar_demux_src2_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_src2_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_src2_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_src2_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_src2_ready),         //          .ready
		.in_data              (cmd_xbar_demux_src2_data),          //          .data
		.out_endofpacket      (width_adapter_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_src_data),            //          .data
		.out_channel          (width_adapter_src_channel),         //          .channel
		.out_valid            (width_adapter_src_valid),           //          .valid
		.out_ready            (width_adapter_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                             // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (106),
		.IN_PKT_RESPONSE_STATUS_L      (105),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (107),
		.OUT_PKT_ADDR_H                (49),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (58),
		.OUT_PKT_BYTE_CNT_L            (56),
		.OUT_PKT_TRANS_COMPRESSED_READ (50),
		.OUT_PKT_BURST_SIZE_H          (64),
		.OUT_PKT_BURST_SIZE_L          (62),
		.OUT_PKT_RESPONSE_STATUS_H     (88),
		.OUT_PKT_RESPONSE_STATUS_L     (87),
		.OUT_PKT_TRANS_EXCLUSIVE       (55),
		.OUT_PKT_BURST_TYPE_H          (66),
		.OUT_PKT_BURST_TYPE_L          (65),
		.OUT_ST_DATA_W                 (89),
		.ST_CHANNEL_W                  (16),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_001 (
		.clk                  (clocks_sys_clk_clk),                    //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (cmd_xbar_demux_001_src2_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_001_src2_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_001_src2_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_001_src2_ready),         //          .ready
		.in_data              (cmd_xbar_demux_001_src2_data),          //          .data
		.out_endofpacket      (width_adapter_001_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_001_src_data),            //          .data
		.out_channel          (width_adapter_001_src_channel),         //          .channel
		.out_valid            (width_adapter_001_src_valid),           //          .valid
		.out_ready            (width_adapter_001_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_001_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (106),
		.IN_PKT_RESPONSE_STATUS_L      (105),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (107),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (49),
		.OUT_PKT_BYTE_CNT_L            (47),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_PKT_BURST_SIZE_H          (55),
		.OUT_PKT_BURST_SIZE_L          (53),
		.OUT_PKT_RESPONSE_STATUS_H     (79),
		.OUT_PKT_RESPONSE_STATUS_L     (78),
		.OUT_PKT_TRANS_EXCLUSIVE       (46),
		.OUT_PKT_BURST_TYPE_H          (57),
		.OUT_PKT_BURST_TYPE_L          (56),
		.OUT_ST_DATA_W                 (80),
		.ST_CHANNEL_W                  (16),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_002 (
		.clk                  (clocks_sys_clk_clk),                    //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (cmd_xbar_demux_001_src9_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_001_src9_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_001_src9_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_001_src9_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_001_src9_ready),         //          .ready
		.in_data              (cmd_xbar_demux_001_src9_data),          //          .data
		.out_endofpacket      (width_adapter_002_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_002_src_data),            //          .data
		.out_channel          (width_adapter_002_src_channel),         //          .channel
		.out_valid            (width_adapter_002_src_valid),           //          .valid
		.out_ready            (width_adapter_002_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_002_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (106),
		.IN_PKT_RESPONSE_STATUS_L      (105),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (107),
		.OUT_PKT_ADDR_H                (49),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (58),
		.OUT_PKT_BYTE_CNT_L            (56),
		.OUT_PKT_TRANS_COMPRESSED_READ (50),
		.OUT_PKT_BURST_SIZE_H          (64),
		.OUT_PKT_BURST_SIZE_L          (62),
		.OUT_PKT_RESPONSE_STATUS_H     (88),
		.OUT_PKT_RESPONSE_STATUS_L     (87),
		.OUT_PKT_TRANS_EXCLUSIVE       (55),
		.OUT_PKT_BURST_TYPE_H          (66),
		.OUT_PKT_BURST_TYPE_L          (65),
		.OUT_ST_DATA_W                 (89),
		.ST_CHANNEL_W                  (16),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_003 (
		.clk                  (clocks_sys_clk_clk),                     //       clk.clk
		.reset                (rst_controller_reset_out_reset),         // clk_reset.reset
		.in_valid             (cmd_xbar_demux_001_src10_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_001_src10_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_001_src10_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_001_src10_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_001_src10_ready),         //          .ready
		.in_data              (cmd_xbar_demux_001_src10_data),          //          .data
		.out_endofpacket      (width_adapter_003_src_endofpacket),      //       src.endofpacket
		.out_data             (width_adapter_003_src_data),             //          .data
		.out_channel          (width_adapter_003_src_channel),          //          .channel
		.out_valid            (width_adapter_003_src_valid),            //          .valid
		.out_ready            (width_adapter_003_src_ready),            //          .ready
		.out_startofpacket    (width_adapter_003_src_startofpacket),    //          .startofpacket
		.in_command_size_data (3'b000)                                  // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (106),
		.IN_PKT_RESPONSE_STATUS_L      (105),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (107),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (49),
		.OUT_PKT_BYTE_CNT_L            (47),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_PKT_BURST_SIZE_H          (55),
		.OUT_PKT_BURST_SIZE_L          (53),
		.OUT_PKT_RESPONSE_STATUS_H     (79),
		.OUT_PKT_RESPONSE_STATUS_L     (78),
		.OUT_PKT_TRANS_EXCLUSIVE       (46),
		.OUT_PKT_BURST_TYPE_H          (57),
		.OUT_PKT_BURST_TYPE_L          (56),
		.OUT_ST_DATA_W                 (80),
		.ST_CHANNEL_W                  (16),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_004 (
		.clk                  (clocks_sys_clk_clk),                     //       clk.clk
		.reset                (rst_controller_reset_out_reset),         // clk_reset.reset
		.in_valid             (cmd_xbar_demux_001_src13_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_001_src13_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_001_src13_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_001_src13_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_001_src13_ready),         //          .ready
		.in_data              (cmd_xbar_demux_001_src13_data),          //          .data
		.out_endofpacket      (width_adapter_004_src_endofpacket),      //       src.endofpacket
		.out_data             (width_adapter_004_src_data),             //          .data
		.out_channel          (width_adapter_004_src_channel),          //          .channel
		.out_valid            (width_adapter_004_src_valid),            //          .valid
		.out_ready            (width_adapter_004_src_ready),            //          .ready
		.out_startofpacket    (width_adapter_004_src_startofpacket),    //          .startofpacket
		.in_command_size_data (3'b000)                                  // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (49),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (58),
		.IN_PKT_BYTE_CNT_L             (56),
		.IN_PKT_TRANS_COMPRESSED_READ  (50),
		.IN_PKT_BURSTWRAP_H            (61),
		.IN_PKT_BURSTWRAP_L            (59),
		.IN_PKT_BURST_SIZE_H           (64),
		.IN_PKT_BURST_SIZE_L           (62),
		.IN_PKT_RESPONSE_STATUS_H      (88),
		.IN_PKT_RESPONSE_STATUS_L      (87),
		.IN_PKT_TRANS_EXCLUSIVE        (55),
		.IN_PKT_BURST_TYPE_H           (66),
		.IN_PKT_BURST_TYPE_L           (65),
		.IN_ST_DATA_W                  (89),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (106),
		.OUT_PKT_RESPONSE_STATUS_L     (105),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (107),
		.ST_CHANNEL_W                  (16),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_005 (
		.clk                  (clocks_sys_clk_clk),                    //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (rsp_xbar_demux_002_src0_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_002_src0_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_002_src0_ready),         //          .ready
		.in_data              (rsp_xbar_demux_002_src0_data),          //          .data
		.out_endofpacket      (width_adapter_005_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_005_src_data),            //          .data
		.out_channel          (width_adapter_005_src_channel),         //          .channel
		.out_valid            (width_adapter_005_src_valid),           //          .valid
		.out_ready            (width_adapter_005_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_005_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (49),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (58),
		.IN_PKT_BYTE_CNT_L             (56),
		.IN_PKT_TRANS_COMPRESSED_READ  (50),
		.IN_PKT_BURSTWRAP_H            (61),
		.IN_PKT_BURSTWRAP_L            (59),
		.IN_PKT_BURST_SIZE_H           (64),
		.IN_PKT_BURST_SIZE_L           (62),
		.IN_PKT_RESPONSE_STATUS_H      (88),
		.IN_PKT_RESPONSE_STATUS_L      (87),
		.IN_PKT_TRANS_EXCLUSIVE        (55),
		.IN_PKT_BURST_TYPE_H           (66),
		.IN_PKT_BURST_TYPE_L           (65),
		.IN_ST_DATA_W                  (89),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (106),
		.OUT_PKT_RESPONSE_STATUS_L     (105),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (107),
		.ST_CHANNEL_W                  (16),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_006 (
		.clk                  (clocks_sys_clk_clk),                    //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (rsp_xbar_demux_002_src1_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_002_src1_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_002_src1_ready),         //          .ready
		.in_data              (rsp_xbar_demux_002_src1_data),          //          .data
		.out_endofpacket      (width_adapter_006_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_006_src_data),            //          .data
		.out_channel          (width_adapter_006_src_channel),         //          .channel
		.out_valid            (width_adapter_006_src_valid),           //          .valid
		.out_ready            (width_adapter_006_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_006_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (49),
		.IN_PKT_BYTE_CNT_L             (47),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (52),
		.IN_PKT_BURSTWRAP_L            (50),
		.IN_PKT_BURST_SIZE_H           (55),
		.IN_PKT_BURST_SIZE_L           (53),
		.IN_PKT_RESPONSE_STATUS_H      (79),
		.IN_PKT_RESPONSE_STATUS_L      (78),
		.IN_PKT_TRANS_EXCLUSIVE        (46),
		.IN_PKT_BURST_TYPE_H           (57),
		.IN_PKT_BURST_TYPE_L           (56),
		.IN_ST_DATA_W                  (80),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (106),
		.OUT_PKT_RESPONSE_STATUS_L     (105),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (107),
		.ST_CHANNEL_W                  (16),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_007 (
		.clk                  (clocks_sys_clk_clk),                    //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (rsp_xbar_demux_009_src0_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_009_src0_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_009_src0_ready),         //          .ready
		.in_data              (rsp_xbar_demux_009_src0_data),          //          .data
		.out_endofpacket      (width_adapter_007_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_007_src_data),            //          .data
		.out_channel          (width_adapter_007_src_channel),         //          .channel
		.out_valid            (width_adapter_007_src_valid),           //          .valid
		.out_ready            (width_adapter_007_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_007_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (49),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (58),
		.IN_PKT_BYTE_CNT_L             (56),
		.IN_PKT_TRANS_COMPRESSED_READ  (50),
		.IN_PKT_BURSTWRAP_H            (61),
		.IN_PKT_BURSTWRAP_L            (59),
		.IN_PKT_BURST_SIZE_H           (64),
		.IN_PKT_BURST_SIZE_L           (62),
		.IN_PKT_RESPONSE_STATUS_H      (88),
		.IN_PKT_RESPONSE_STATUS_L      (87),
		.IN_PKT_TRANS_EXCLUSIVE        (55),
		.IN_PKT_BURST_TYPE_H           (66),
		.IN_PKT_BURST_TYPE_L           (65),
		.IN_ST_DATA_W                  (89),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (106),
		.OUT_PKT_RESPONSE_STATUS_L     (105),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (107),
		.ST_CHANNEL_W                  (16),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_008 (
		.clk                  (clocks_sys_clk_clk),                    //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (rsp_xbar_demux_010_src0_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_010_src0_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_010_src0_ready),         //          .ready
		.in_data              (rsp_xbar_demux_010_src0_data),          //          .data
		.out_endofpacket      (width_adapter_008_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_008_src_data),            //          .data
		.out_channel          (width_adapter_008_src_channel),         //          .channel
		.out_valid            (width_adapter_008_src_valid),           //          .valid
		.out_ready            (width_adapter_008_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_008_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (49),
		.IN_PKT_BYTE_CNT_L             (47),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (52),
		.IN_PKT_BURSTWRAP_L            (50),
		.IN_PKT_BURST_SIZE_H           (55),
		.IN_PKT_BURST_SIZE_L           (53),
		.IN_PKT_RESPONSE_STATUS_H      (79),
		.IN_PKT_RESPONSE_STATUS_L      (78),
		.IN_PKT_TRANS_EXCLUSIVE        (46),
		.IN_PKT_BURST_TYPE_H           (57),
		.IN_PKT_BURST_TYPE_L           (56),
		.IN_ST_DATA_W                  (80),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (106),
		.OUT_PKT_RESPONSE_STATUS_L     (105),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (107),
		.ST_CHANNEL_W                  (16),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_009 (
		.clk                  (clocks_sys_clk_clk),                    //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (rsp_xbar_demux_013_src0_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_013_src0_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_013_src0_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_013_src0_ready),         //          .ready
		.in_data              (rsp_xbar_demux_013_src0_data),          //          .data
		.out_endofpacket      (width_adapter_009_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_009_src_data),            //          .data
		.out_channel          (width_adapter_009_src_channel),         //          .channel
		.out_valid            (width_adapter_009_src_valid),           //          .valid
		.out_ready            (width_adapter_009_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_009_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	nios_system_irq_mapper irq_mapper (
		.clk           (clocks_sys_clk_clk),             //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.sender_irq    (nios2_qsys_0_d_irq_irq)          //    sender.irq
	);

endmodule
